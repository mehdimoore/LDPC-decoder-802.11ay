always @(posedge clk)begin
if (chk_n_output_valid[0] & active_cols[0]) begin
case (curr_layer)
    0:begin 
        eta_sum[0][40]  = eta_sum_out_tmp[0][0];
        eta_sum[0][41]  = eta_sum_out_tmp[0][1];
        eta_sum[0][0]  = eta_sum_out_tmp[0][2];
        eta_sum[0][1]  = eta_sum_out_tmp[0][3];
        eta_sum[0][2]  = eta_sum_out_tmp[0][4];
        eta_sum[0][3]  = eta_sum_out_tmp[0][5];
        eta_sum[0][4]  = eta_sum_out_tmp[0][6];
        eta_sum[0][5]  = eta_sum_out_tmp[0][7];
        eta_sum[0][6]  = eta_sum_out_tmp[0][8];
        eta_sum[0][7]  = eta_sum_out_tmp[0][9];
        eta_sum[0][8]  = eta_sum_out_tmp[0][10];
        eta_sum[0][9]  = eta_sum_out_tmp[0][11];
        eta_sum[0][10]  = eta_sum_out_tmp[0][12];
        eta_sum[0][11]  = eta_sum_out_tmp[0][13];
        eta_sum[0][12]  = eta_sum_out_tmp[0][14];
        eta_sum[0][13]  = eta_sum_out_tmp[0][15];
        eta_sum[0][14]  = eta_sum_out_tmp[0][16];
        eta_sum[0][15]  = eta_sum_out_tmp[0][17];
        eta_sum[0][16]  = eta_sum_out_tmp[0][18];
        eta_sum[0][17]  = eta_sum_out_tmp[0][19];
        eta_sum[0][18]  = eta_sum_out_tmp[0][20];
        eta_sum[0][19]  = eta_sum_out_tmp[0][21];
        eta_sum[0][20]  = eta_sum_out_tmp[0][22];
        eta_sum[0][21]  = eta_sum_out_tmp[0][23];
        eta_sum[0][22]  = eta_sum_out_tmp[0][24];
        eta_sum[0][23]  = eta_sum_out_tmp[0][25];
        eta_sum[0][24]  = eta_sum_out_tmp[0][26];
        eta_sum[0][25]  = eta_sum_out_tmp[0][27];
        eta_sum[0][26]  = eta_sum_out_tmp[0][28];
        eta_sum[0][27]  = eta_sum_out_tmp[0][29];
        eta_sum[0][28]  = eta_sum_out_tmp[0][30];
        eta_sum[0][29]  = eta_sum_out_tmp[0][31];
        eta_sum[0][30]  = eta_sum_out_tmp[0][32];
        eta_sum[0][31]  = eta_sum_out_tmp[0][33];
        eta_sum[0][32]  = eta_sum_out_tmp[0][34];
        eta_sum[0][33]  = eta_sum_out_tmp[0][35];
        eta_sum[0][34]  = eta_sum_out_tmp[0][36];
        eta_sum[0][35]  = eta_sum_out_tmp[0][37];
        eta_sum[0][36]  = eta_sum_out_tmp[0][38];
        eta_sum[0][37]  = eta_sum_out_tmp[0][39];
        eta_sum[0][38]  = eta_sum_out_tmp[0][40];
        eta_sum[0][39]  = eta_sum_out_tmp[0][41];
    end
 
    1:begin 
        eta_sum[0][34]  = eta_sum_out_tmp[0][0];
        eta_sum[0][35]  = eta_sum_out_tmp[0][1];
        eta_sum[0][36]  = eta_sum_out_tmp[0][2];
        eta_sum[0][37]  = eta_sum_out_tmp[0][3];
        eta_sum[0][38]  = eta_sum_out_tmp[0][4];
        eta_sum[0][39]  = eta_sum_out_tmp[0][5];
        eta_sum[0][40]  = eta_sum_out_tmp[0][6];
        eta_sum[0][41]  = eta_sum_out_tmp[0][7];
        eta_sum[0][0]  = eta_sum_out_tmp[0][8];
        eta_sum[0][1]  = eta_sum_out_tmp[0][9];
        eta_sum[0][2]  = eta_sum_out_tmp[0][10];
        eta_sum[0][3]  = eta_sum_out_tmp[0][11];
        eta_sum[0][4]  = eta_sum_out_tmp[0][12];
        eta_sum[0][5]  = eta_sum_out_tmp[0][13];
        eta_sum[0][6]  = eta_sum_out_tmp[0][14];
        eta_sum[0][7]  = eta_sum_out_tmp[0][15];
        eta_sum[0][8]  = eta_sum_out_tmp[0][16];
        eta_sum[0][9]  = eta_sum_out_tmp[0][17];
        eta_sum[0][10]  = eta_sum_out_tmp[0][18];
        eta_sum[0][11]  = eta_sum_out_tmp[0][19];
        eta_sum[0][12]  = eta_sum_out_tmp[0][20];
        eta_sum[0][13]  = eta_sum_out_tmp[0][21];
        eta_sum[0][14]  = eta_sum_out_tmp[0][22];
        eta_sum[0][15]  = eta_sum_out_tmp[0][23];
        eta_sum[0][16]  = eta_sum_out_tmp[0][24];
        eta_sum[0][17]  = eta_sum_out_tmp[0][25];
        eta_sum[0][18]  = eta_sum_out_tmp[0][26];
        eta_sum[0][19]  = eta_sum_out_tmp[0][27];
        eta_sum[0][20]  = eta_sum_out_tmp[0][28];
        eta_sum[0][21]  = eta_sum_out_tmp[0][29];
        eta_sum[0][22]  = eta_sum_out_tmp[0][30];
        eta_sum[0][23]  = eta_sum_out_tmp[0][31];
        eta_sum[0][24]  = eta_sum_out_tmp[0][32];
        eta_sum[0][25]  = eta_sum_out_tmp[0][33];
        eta_sum[0][26]  = eta_sum_out_tmp[0][34];
        eta_sum[0][27]  = eta_sum_out_tmp[0][35];
        eta_sum[0][28]  = eta_sum_out_tmp[0][36];
        eta_sum[0][29]  = eta_sum_out_tmp[0][37];
        eta_sum[0][30]  = eta_sum_out_tmp[0][38];
        eta_sum[0][31]  = eta_sum_out_tmp[0][39];
        eta_sum[0][32]  = eta_sum_out_tmp[0][40];
        eta_sum[0][33]  = eta_sum_out_tmp[0][41];
    end
 
    2:begin 
        eta_sum[0][0]  = eta_sum_out_tmp[0][0];
        eta_sum[0][1]  = eta_sum_out_tmp[0][1];
        eta_sum[0][2]  = eta_sum_out_tmp[0][2];
        eta_sum[0][3]  = eta_sum_out_tmp[0][3];
        eta_sum[0][4]  = eta_sum_out_tmp[0][4];
        eta_sum[0][5]  = eta_sum_out_tmp[0][5];
        eta_sum[0][6]  = eta_sum_out_tmp[0][6];
        eta_sum[0][7]  = eta_sum_out_tmp[0][7];
        eta_sum[0][8]  = eta_sum_out_tmp[0][8];
        eta_sum[0][9]  = eta_sum_out_tmp[0][9];
        eta_sum[0][10]  = eta_sum_out_tmp[0][10];
        eta_sum[0][11]  = eta_sum_out_tmp[0][11];
        eta_sum[0][12]  = eta_sum_out_tmp[0][12];
        eta_sum[0][13]  = eta_sum_out_tmp[0][13];
        eta_sum[0][14]  = eta_sum_out_tmp[0][14];
        eta_sum[0][15]  = eta_sum_out_tmp[0][15];
        eta_sum[0][16]  = eta_sum_out_tmp[0][16];
        eta_sum[0][17]  = eta_sum_out_tmp[0][17];
        eta_sum[0][18]  = eta_sum_out_tmp[0][18];
        eta_sum[0][19]  = eta_sum_out_tmp[0][19];
        eta_sum[0][20]  = eta_sum_out_tmp[0][20];
        eta_sum[0][21]  = eta_sum_out_tmp[0][21];
        eta_sum[0][22]  = eta_sum_out_tmp[0][22];
        eta_sum[0][23]  = eta_sum_out_tmp[0][23];
        eta_sum[0][24]  = eta_sum_out_tmp[0][24];
        eta_sum[0][25]  = eta_sum_out_tmp[0][25];
        eta_sum[0][26]  = eta_sum_out_tmp[0][26];
        eta_sum[0][27]  = eta_sum_out_tmp[0][27];
        eta_sum[0][28]  = eta_sum_out_tmp[0][28];
        eta_sum[0][29]  = eta_sum_out_tmp[0][29];
        eta_sum[0][30]  = eta_sum_out_tmp[0][30];
        eta_sum[0][31]  = eta_sum_out_tmp[0][31];
        eta_sum[0][32]  = eta_sum_out_tmp[0][32];
        eta_sum[0][33]  = eta_sum_out_tmp[0][33];
        eta_sum[0][34]  = eta_sum_out_tmp[0][34];
        eta_sum[0][35]  = eta_sum_out_tmp[0][35];
        eta_sum[0][36]  = eta_sum_out_tmp[0][36];
        eta_sum[0][37]  = eta_sum_out_tmp[0][37];
        eta_sum[0][38]  = eta_sum_out_tmp[0][38];
        eta_sum[0][39]  = eta_sum_out_tmp[0][39];
        eta_sum[0][40]  = eta_sum_out_tmp[0][40];
        eta_sum[0][41]  = eta_sum_out_tmp[0][41];
    end
 
    3:begin 
        eta_sum[0][0]  = eta_sum_out_tmp[0][0];
        eta_sum[0][1]  = eta_sum_out_tmp[0][1];
        eta_sum[0][2]  = eta_sum_out_tmp[0][2];
        eta_sum[0][3]  = eta_sum_out_tmp[0][3];
        eta_sum[0][4]  = eta_sum_out_tmp[0][4];
        eta_sum[0][5]  = eta_sum_out_tmp[0][5];
        eta_sum[0][6]  = eta_sum_out_tmp[0][6];
        eta_sum[0][7]  = eta_sum_out_tmp[0][7];
        eta_sum[0][8]  = eta_sum_out_tmp[0][8];
        eta_sum[0][9]  = eta_sum_out_tmp[0][9];
        eta_sum[0][10]  = eta_sum_out_tmp[0][10];
        eta_sum[0][11]  = eta_sum_out_tmp[0][11];
        eta_sum[0][12]  = eta_sum_out_tmp[0][12];
        eta_sum[0][13]  = eta_sum_out_tmp[0][13];
        eta_sum[0][14]  = eta_sum_out_tmp[0][14];
        eta_sum[0][15]  = eta_sum_out_tmp[0][15];
        eta_sum[0][16]  = eta_sum_out_tmp[0][16];
        eta_sum[0][17]  = eta_sum_out_tmp[0][17];
        eta_sum[0][18]  = eta_sum_out_tmp[0][18];
        eta_sum[0][19]  = eta_sum_out_tmp[0][19];
        eta_sum[0][20]  = eta_sum_out_tmp[0][20];
        eta_sum[0][21]  = eta_sum_out_tmp[0][21];
        eta_sum[0][22]  = eta_sum_out_tmp[0][22];
        eta_sum[0][23]  = eta_sum_out_tmp[0][23];
        eta_sum[0][24]  = eta_sum_out_tmp[0][24];
        eta_sum[0][25]  = eta_sum_out_tmp[0][25];
        eta_sum[0][26]  = eta_sum_out_tmp[0][26];
        eta_sum[0][27]  = eta_sum_out_tmp[0][27];
        eta_sum[0][28]  = eta_sum_out_tmp[0][28];
        eta_sum[0][29]  = eta_sum_out_tmp[0][29];
        eta_sum[0][30]  = eta_sum_out_tmp[0][30];
        eta_sum[0][31]  = eta_sum_out_tmp[0][31];
        eta_sum[0][32]  = eta_sum_out_tmp[0][32];
        eta_sum[0][33]  = eta_sum_out_tmp[0][33];
        eta_sum[0][34]  = eta_sum_out_tmp[0][34];
        eta_sum[0][35]  = eta_sum_out_tmp[0][35];
        eta_sum[0][36]  = eta_sum_out_tmp[0][36];
        eta_sum[0][37]  = eta_sum_out_tmp[0][37];
        eta_sum[0][38]  = eta_sum_out_tmp[0][38];
        eta_sum[0][39]  = eta_sum_out_tmp[0][39];
        eta_sum[0][40]  = eta_sum_out_tmp[0][40];
        eta_sum[0][41]  = eta_sum_out_tmp[0][41];
    end
 
    4:begin 
        eta_sum[0][35]  = eta_sum_out_tmp[0][0];
        eta_sum[0][36]  = eta_sum_out_tmp[0][1];
        eta_sum[0][37]  = eta_sum_out_tmp[0][2];
        eta_sum[0][38]  = eta_sum_out_tmp[0][3];
        eta_sum[0][39]  = eta_sum_out_tmp[0][4];
        eta_sum[0][40]  = eta_sum_out_tmp[0][5];
        eta_sum[0][41]  = eta_sum_out_tmp[0][6];
        eta_sum[0][0]  = eta_sum_out_tmp[0][7];
        eta_sum[0][1]  = eta_sum_out_tmp[0][8];
        eta_sum[0][2]  = eta_sum_out_tmp[0][9];
        eta_sum[0][3]  = eta_sum_out_tmp[0][10];
        eta_sum[0][4]  = eta_sum_out_tmp[0][11];
        eta_sum[0][5]  = eta_sum_out_tmp[0][12];
        eta_sum[0][6]  = eta_sum_out_tmp[0][13];
        eta_sum[0][7]  = eta_sum_out_tmp[0][14];
        eta_sum[0][8]  = eta_sum_out_tmp[0][15];
        eta_sum[0][9]  = eta_sum_out_tmp[0][16];
        eta_sum[0][10]  = eta_sum_out_tmp[0][17];
        eta_sum[0][11]  = eta_sum_out_tmp[0][18];
        eta_sum[0][12]  = eta_sum_out_tmp[0][19];
        eta_sum[0][13]  = eta_sum_out_tmp[0][20];
        eta_sum[0][14]  = eta_sum_out_tmp[0][21];
        eta_sum[0][15]  = eta_sum_out_tmp[0][22];
        eta_sum[0][16]  = eta_sum_out_tmp[0][23];
        eta_sum[0][17]  = eta_sum_out_tmp[0][24];
        eta_sum[0][18]  = eta_sum_out_tmp[0][25];
        eta_sum[0][19]  = eta_sum_out_tmp[0][26];
        eta_sum[0][20]  = eta_sum_out_tmp[0][27];
        eta_sum[0][21]  = eta_sum_out_tmp[0][28];
        eta_sum[0][22]  = eta_sum_out_tmp[0][29];
        eta_sum[0][23]  = eta_sum_out_tmp[0][30];
        eta_sum[0][24]  = eta_sum_out_tmp[0][31];
        eta_sum[0][25]  = eta_sum_out_tmp[0][32];
        eta_sum[0][26]  = eta_sum_out_tmp[0][33];
        eta_sum[0][27]  = eta_sum_out_tmp[0][34];
        eta_sum[0][28]  = eta_sum_out_tmp[0][35];
        eta_sum[0][29]  = eta_sum_out_tmp[0][36];
        eta_sum[0][30]  = eta_sum_out_tmp[0][37];
        eta_sum[0][31]  = eta_sum_out_tmp[0][38];
        eta_sum[0][32]  = eta_sum_out_tmp[0][39];
        eta_sum[0][33]  = eta_sum_out_tmp[0][40];
        eta_sum[0][34]  = eta_sum_out_tmp[0][41];
    end
 
    5:begin 
        eta_sum[0][29]  = eta_sum_out_tmp[0][0];
        eta_sum[0][30]  = eta_sum_out_tmp[0][1];
        eta_sum[0][31]  = eta_sum_out_tmp[0][2];
        eta_sum[0][32]  = eta_sum_out_tmp[0][3];
        eta_sum[0][33]  = eta_sum_out_tmp[0][4];
        eta_sum[0][34]  = eta_sum_out_tmp[0][5];
        eta_sum[0][35]  = eta_sum_out_tmp[0][6];
        eta_sum[0][36]  = eta_sum_out_tmp[0][7];
        eta_sum[0][37]  = eta_sum_out_tmp[0][8];
        eta_sum[0][38]  = eta_sum_out_tmp[0][9];
        eta_sum[0][39]  = eta_sum_out_tmp[0][10];
        eta_sum[0][40]  = eta_sum_out_tmp[0][11];
        eta_sum[0][41]  = eta_sum_out_tmp[0][12];
        eta_sum[0][0]  = eta_sum_out_tmp[0][13];
        eta_sum[0][1]  = eta_sum_out_tmp[0][14];
        eta_sum[0][2]  = eta_sum_out_tmp[0][15];
        eta_sum[0][3]  = eta_sum_out_tmp[0][16];
        eta_sum[0][4]  = eta_sum_out_tmp[0][17];
        eta_sum[0][5]  = eta_sum_out_tmp[0][18];
        eta_sum[0][6]  = eta_sum_out_tmp[0][19];
        eta_sum[0][7]  = eta_sum_out_tmp[0][20];
        eta_sum[0][8]  = eta_sum_out_tmp[0][21];
        eta_sum[0][9]  = eta_sum_out_tmp[0][22];
        eta_sum[0][10]  = eta_sum_out_tmp[0][23];
        eta_sum[0][11]  = eta_sum_out_tmp[0][24];
        eta_sum[0][12]  = eta_sum_out_tmp[0][25];
        eta_sum[0][13]  = eta_sum_out_tmp[0][26];
        eta_sum[0][14]  = eta_sum_out_tmp[0][27];
        eta_sum[0][15]  = eta_sum_out_tmp[0][28];
        eta_sum[0][16]  = eta_sum_out_tmp[0][29];
        eta_sum[0][17]  = eta_sum_out_tmp[0][30];
        eta_sum[0][18]  = eta_sum_out_tmp[0][31];
        eta_sum[0][19]  = eta_sum_out_tmp[0][32];
        eta_sum[0][20]  = eta_sum_out_tmp[0][33];
        eta_sum[0][21]  = eta_sum_out_tmp[0][34];
        eta_sum[0][22]  = eta_sum_out_tmp[0][35];
        eta_sum[0][23]  = eta_sum_out_tmp[0][36];
        eta_sum[0][24]  = eta_sum_out_tmp[0][37];
        eta_sum[0][25]  = eta_sum_out_tmp[0][38];
        eta_sum[0][26]  = eta_sum_out_tmp[0][39];
        eta_sum[0][27]  = eta_sum_out_tmp[0][40];
        eta_sum[0][28]  = eta_sum_out_tmp[0][41];
    end
 
    6:begin 
        eta_sum[0][0]  = eta_sum_out_tmp[0][0];
        eta_sum[0][1]  = eta_sum_out_tmp[0][1];
        eta_sum[0][2]  = eta_sum_out_tmp[0][2];
        eta_sum[0][3]  = eta_sum_out_tmp[0][3];
        eta_sum[0][4]  = eta_sum_out_tmp[0][4];
        eta_sum[0][5]  = eta_sum_out_tmp[0][5];
        eta_sum[0][6]  = eta_sum_out_tmp[0][6];
        eta_sum[0][7]  = eta_sum_out_tmp[0][7];
        eta_sum[0][8]  = eta_sum_out_tmp[0][8];
        eta_sum[0][9]  = eta_sum_out_tmp[0][9];
        eta_sum[0][10]  = eta_sum_out_tmp[0][10];
        eta_sum[0][11]  = eta_sum_out_tmp[0][11];
        eta_sum[0][12]  = eta_sum_out_tmp[0][12];
        eta_sum[0][13]  = eta_sum_out_tmp[0][13];
        eta_sum[0][14]  = eta_sum_out_tmp[0][14];
        eta_sum[0][15]  = eta_sum_out_tmp[0][15];
        eta_sum[0][16]  = eta_sum_out_tmp[0][16];
        eta_sum[0][17]  = eta_sum_out_tmp[0][17];
        eta_sum[0][18]  = eta_sum_out_tmp[0][18];
        eta_sum[0][19]  = eta_sum_out_tmp[0][19];
        eta_sum[0][20]  = eta_sum_out_tmp[0][20];
        eta_sum[0][21]  = eta_sum_out_tmp[0][21];
        eta_sum[0][22]  = eta_sum_out_tmp[0][22];
        eta_sum[0][23]  = eta_sum_out_tmp[0][23];
        eta_sum[0][24]  = eta_sum_out_tmp[0][24];
        eta_sum[0][25]  = eta_sum_out_tmp[0][25];
        eta_sum[0][26]  = eta_sum_out_tmp[0][26];
        eta_sum[0][27]  = eta_sum_out_tmp[0][27];
        eta_sum[0][28]  = eta_sum_out_tmp[0][28];
        eta_sum[0][29]  = eta_sum_out_tmp[0][29];
        eta_sum[0][30]  = eta_sum_out_tmp[0][30];
        eta_sum[0][31]  = eta_sum_out_tmp[0][31];
        eta_sum[0][32]  = eta_sum_out_tmp[0][32];
        eta_sum[0][33]  = eta_sum_out_tmp[0][33];
        eta_sum[0][34]  = eta_sum_out_tmp[0][34];
        eta_sum[0][35]  = eta_sum_out_tmp[0][35];
        eta_sum[0][36]  = eta_sum_out_tmp[0][36];
        eta_sum[0][37]  = eta_sum_out_tmp[0][37];
        eta_sum[0][38]  = eta_sum_out_tmp[0][38];
        eta_sum[0][39]  = eta_sum_out_tmp[0][39];
        eta_sum[0][40]  = eta_sum_out_tmp[0][40];
        eta_sum[0][41]  = eta_sum_out_tmp[0][41];
    end
 
    7:begin 
        eta_sum[0][0]  = eta_sum_out_tmp[0][0];
        eta_sum[0][1]  = eta_sum_out_tmp[0][1];
        eta_sum[0][2]  = eta_sum_out_tmp[0][2];
        eta_sum[0][3]  = eta_sum_out_tmp[0][3];
        eta_sum[0][4]  = eta_sum_out_tmp[0][4];
        eta_sum[0][5]  = eta_sum_out_tmp[0][5];
        eta_sum[0][6]  = eta_sum_out_tmp[0][6];
        eta_sum[0][7]  = eta_sum_out_tmp[0][7];
        eta_sum[0][8]  = eta_sum_out_tmp[0][8];
        eta_sum[0][9]  = eta_sum_out_tmp[0][9];
        eta_sum[0][10]  = eta_sum_out_tmp[0][10];
        eta_sum[0][11]  = eta_sum_out_tmp[0][11];
        eta_sum[0][12]  = eta_sum_out_tmp[0][12];
        eta_sum[0][13]  = eta_sum_out_tmp[0][13];
        eta_sum[0][14]  = eta_sum_out_tmp[0][14];
        eta_sum[0][15]  = eta_sum_out_tmp[0][15];
        eta_sum[0][16]  = eta_sum_out_tmp[0][16];
        eta_sum[0][17]  = eta_sum_out_tmp[0][17];
        eta_sum[0][18]  = eta_sum_out_tmp[0][18];
        eta_sum[0][19]  = eta_sum_out_tmp[0][19];
        eta_sum[0][20]  = eta_sum_out_tmp[0][20];
        eta_sum[0][21]  = eta_sum_out_tmp[0][21];
        eta_sum[0][22]  = eta_sum_out_tmp[0][22];
        eta_sum[0][23]  = eta_sum_out_tmp[0][23];
        eta_sum[0][24]  = eta_sum_out_tmp[0][24];
        eta_sum[0][25]  = eta_sum_out_tmp[0][25];
        eta_sum[0][26]  = eta_sum_out_tmp[0][26];
        eta_sum[0][27]  = eta_sum_out_tmp[0][27];
        eta_sum[0][28]  = eta_sum_out_tmp[0][28];
        eta_sum[0][29]  = eta_sum_out_tmp[0][29];
        eta_sum[0][30]  = eta_sum_out_tmp[0][30];
        eta_sum[0][31]  = eta_sum_out_tmp[0][31];
        eta_sum[0][32]  = eta_sum_out_tmp[0][32];
        eta_sum[0][33]  = eta_sum_out_tmp[0][33];
        eta_sum[0][34]  = eta_sum_out_tmp[0][34];
        eta_sum[0][35]  = eta_sum_out_tmp[0][35];
        eta_sum[0][36]  = eta_sum_out_tmp[0][36];
        eta_sum[0][37]  = eta_sum_out_tmp[0][37];
        eta_sum[0][38]  = eta_sum_out_tmp[0][38];
        eta_sum[0][39]  = eta_sum_out_tmp[0][39];
        eta_sum[0][40]  = eta_sum_out_tmp[0][40];
        eta_sum[0][41]  = eta_sum_out_tmp[0][41];
    end
endcase
end

if (chk_n_output_valid[0] & active_cols[1]) begin
case (curr_layer)
    0:begin 
        eta_sum[1][0]  = eta_sum_out_tmp[1][0];
        eta_sum[1][1]  = eta_sum_out_tmp[1][1];
        eta_sum[1][2]  = eta_sum_out_tmp[1][2];
        eta_sum[1][3]  = eta_sum_out_tmp[1][3];
        eta_sum[1][4]  = eta_sum_out_tmp[1][4];
        eta_sum[1][5]  = eta_sum_out_tmp[1][5];
        eta_sum[1][6]  = eta_sum_out_tmp[1][6];
        eta_sum[1][7]  = eta_sum_out_tmp[1][7];
        eta_sum[1][8]  = eta_sum_out_tmp[1][8];
        eta_sum[1][9]  = eta_sum_out_tmp[1][9];
        eta_sum[1][10]  = eta_sum_out_tmp[1][10];
        eta_sum[1][11]  = eta_sum_out_tmp[1][11];
        eta_sum[1][12]  = eta_sum_out_tmp[1][12];
        eta_sum[1][13]  = eta_sum_out_tmp[1][13];
        eta_sum[1][14]  = eta_sum_out_tmp[1][14];
        eta_sum[1][15]  = eta_sum_out_tmp[1][15];
        eta_sum[1][16]  = eta_sum_out_tmp[1][16];
        eta_sum[1][17]  = eta_sum_out_tmp[1][17];
        eta_sum[1][18]  = eta_sum_out_tmp[1][18];
        eta_sum[1][19]  = eta_sum_out_tmp[1][19];
        eta_sum[1][20]  = eta_sum_out_tmp[1][20];
        eta_sum[1][21]  = eta_sum_out_tmp[1][21];
        eta_sum[1][22]  = eta_sum_out_tmp[1][22];
        eta_sum[1][23]  = eta_sum_out_tmp[1][23];
        eta_sum[1][24]  = eta_sum_out_tmp[1][24];
        eta_sum[1][25]  = eta_sum_out_tmp[1][25];
        eta_sum[1][26]  = eta_sum_out_tmp[1][26];
        eta_sum[1][27]  = eta_sum_out_tmp[1][27];
        eta_sum[1][28]  = eta_sum_out_tmp[1][28];
        eta_sum[1][29]  = eta_sum_out_tmp[1][29];
        eta_sum[1][30]  = eta_sum_out_tmp[1][30];
        eta_sum[1][31]  = eta_sum_out_tmp[1][31];
        eta_sum[1][32]  = eta_sum_out_tmp[1][32];
        eta_sum[1][33]  = eta_sum_out_tmp[1][33];
        eta_sum[1][34]  = eta_sum_out_tmp[1][34];
        eta_sum[1][35]  = eta_sum_out_tmp[1][35];
        eta_sum[1][36]  = eta_sum_out_tmp[1][36];
        eta_sum[1][37]  = eta_sum_out_tmp[1][37];
        eta_sum[1][38]  = eta_sum_out_tmp[1][38];
        eta_sum[1][39]  = eta_sum_out_tmp[1][39];
        eta_sum[1][40]  = eta_sum_out_tmp[1][40];
        eta_sum[1][41]  = eta_sum_out_tmp[1][41];
    end
 
    1:begin 
        eta_sum[1][0]  = eta_sum_out_tmp[1][0];
        eta_sum[1][1]  = eta_sum_out_tmp[1][1];
        eta_sum[1][2]  = eta_sum_out_tmp[1][2];
        eta_sum[1][3]  = eta_sum_out_tmp[1][3];
        eta_sum[1][4]  = eta_sum_out_tmp[1][4];
        eta_sum[1][5]  = eta_sum_out_tmp[1][5];
        eta_sum[1][6]  = eta_sum_out_tmp[1][6];
        eta_sum[1][7]  = eta_sum_out_tmp[1][7];
        eta_sum[1][8]  = eta_sum_out_tmp[1][8];
        eta_sum[1][9]  = eta_sum_out_tmp[1][9];
        eta_sum[1][10]  = eta_sum_out_tmp[1][10];
        eta_sum[1][11]  = eta_sum_out_tmp[1][11];
        eta_sum[1][12]  = eta_sum_out_tmp[1][12];
        eta_sum[1][13]  = eta_sum_out_tmp[1][13];
        eta_sum[1][14]  = eta_sum_out_tmp[1][14];
        eta_sum[1][15]  = eta_sum_out_tmp[1][15];
        eta_sum[1][16]  = eta_sum_out_tmp[1][16];
        eta_sum[1][17]  = eta_sum_out_tmp[1][17];
        eta_sum[1][18]  = eta_sum_out_tmp[1][18];
        eta_sum[1][19]  = eta_sum_out_tmp[1][19];
        eta_sum[1][20]  = eta_sum_out_tmp[1][20];
        eta_sum[1][21]  = eta_sum_out_tmp[1][21];
        eta_sum[1][22]  = eta_sum_out_tmp[1][22];
        eta_sum[1][23]  = eta_sum_out_tmp[1][23];
        eta_sum[1][24]  = eta_sum_out_tmp[1][24];
        eta_sum[1][25]  = eta_sum_out_tmp[1][25];
        eta_sum[1][26]  = eta_sum_out_tmp[1][26];
        eta_sum[1][27]  = eta_sum_out_tmp[1][27];
        eta_sum[1][28]  = eta_sum_out_tmp[1][28];
        eta_sum[1][29]  = eta_sum_out_tmp[1][29];
        eta_sum[1][30]  = eta_sum_out_tmp[1][30];
        eta_sum[1][31]  = eta_sum_out_tmp[1][31];
        eta_sum[1][32]  = eta_sum_out_tmp[1][32];
        eta_sum[1][33]  = eta_sum_out_tmp[1][33];
        eta_sum[1][34]  = eta_sum_out_tmp[1][34];
        eta_sum[1][35]  = eta_sum_out_tmp[1][35];
        eta_sum[1][36]  = eta_sum_out_tmp[1][36];
        eta_sum[1][37]  = eta_sum_out_tmp[1][37];
        eta_sum[1][38]  = eta_sum_out_tmp[1][38];
        eta_sum[1][39]  = eta_sum_out_tmp[1][39];
        eta_sum[1][40]  = eta_sum_out_tmp[1][40];
        eta_sum[1][41]  = eta_sum_out_tmp[1][41];
    end
 
    2:begin 
        eta_sum[1][36]  = eta_sum_out_tmp[1][0];
        eta_sum[1][37]  = eta_sum_out_tmp[1][1];
        eta_sum[1][38]  = eta_sum_out_tmp[1][2];
        eta_sum[1][39]  = eta_sum_out_tmp[1][3];
        eta_sum[1][40]  = eta_sum_out_tmp[1][4];
        eta_sum[1][41]  = eta_sum_out_tmp[1][5];
        eta_sum[1][0]  = eta_sum_out_tmp[1][6];
        eta_sum[1][1]  = eta_sum_out_tmp[1][7];
        eta_sum[1][2]  = eta_sum_out_tmp[1][8];
        eta_sum[1][3]  = eta_sum_out_tmp[1][9];
        eta_sum[1][4]  = eta_sum_out_tmp[1][10];
        eta_sum[1][5]  = eta_sum_out_tmp[1][11];
        eta_sum[1][6]  = eta_sum_out_tmp[1][12];
        eta_sum[1][7]  = eta_sum_out_tmp[1][13];
        eta_sum[1][8]  = eta_sum_out_tmp[1][14];
        eta_sum[1][9]  = eta_sum_out_tmp[1][15];
        eta_sum[1][10]  = eta_sum_out_tmp[1][16];
        eta_sum[1][11]  = eta_sum_out_tmp[1][17];
        eta_sum[1][12]  = eta_sum_out_tmp[1][18];
        eta_sum[1][13]  = eta_sum_out_tmp[1][19];
        eta_sum[1][14]  = eta_sum_out_tmp[1][20];
        eta_sum[1][15]  = eta_sum_out_tmp[1][21];
        eta_sum[1][16]  = eta_sum_out_tmp[1][22];
        eta_sum[1][17]  = eta_sum_out_tmp[1][23];
        eta_sum[1][18]  = eta_sum_out_tmp[1][24];
        eta_sum[1][19]  = eta_sum_out_tmp[1][25];
        eta_sum[1][20]  = eta_sum_out_tmp[1][26];
        eta_sum[1][21]  = eta_sum_out_tmp[1][27];
        eta_sum[1][22]  = eta_sum_out_tmp[1][28];
        eta_sum[1][23]  = eta_sum_out_tmp[1][29];
        eta_sum[1][24]  = eta_sum_out_tmp[1][30];
        eta_sum[1][25]  = eta_sum_out_tmp[1][31];
        eta_sum[1][26]  = eta_sum_out_tmp[1][32];
        eta_sum[1][27]  = eta_sum_out_tmp[1][33];
        eta_sum[1][28]  = eta_sum_out_tmp[1][34];
        eta_sum[1][29]  = eta_sum_out_tmp[1][35];
        eta_sum[1][30]  = eta_sum_out_tmp[1][36];
        eta_sum[1][31]  = eta_sum_out_tmp[1][37];
        eta_sum[1][32]  = eta_sum_out_tmp[1][38];
        eta_sum[1][33]  = eta_sum_out_tmp[1][39];
        eta_sum[1][34]  = eta_sum_out_tmp[1][40];
        eta_sum[1][35]  = eta_sum_out_tmp[1][41];
    end
 
    3:begin 
        eta_sum[1][27]  = eta_sum_out_tmp[1][0];
        eta_sum[1][28]  = eta_sum_out_tmp[1][1];
        eta_sum[1][29]  = eta_sum_out_tmp[1][2];
        eta_sum[1][30]  = eta_sum_out_tmp[1][3];
        eta_sum[1][31]  = eta_sum_out_tmp[1][4];
        eta_sum[1][32]  = eta_sum_out_tmp[1][5];
        eta_sum[1][33]  = eta_sum_out_tmp[1][6];
        eta_sum[1][34]  = eta_sum_out_tmp[1][7];
        eta_sum[1][35]  = eta_sum_out_tmp[1][8];
        eta_sum[1][36]  = eta_sum_out_tmp[1][9];
        eta_sum[1][37]  = eta_sum_out_tmp[1][10];
        eta_sum[1][38]  = eta_sum_out_tmp[1][11];
        eta_sum[1][39]  = eta_sum_out_tmp[1][12];
        eta_sum[1][40]  = eta_sum_out_tmp[1][13];
        eta_sum[1][41]  = eta_sum_out_tmp[1][14];
        eta_sum[1][0]  = eta_sum_out_tmp[1][15];
        eta_sum[1][1]  = eta_sum_out_tmp[1][16];
        eta_sum[1][2]  = eta_sum_out_tmp[1][17];
        eta_sum[1][3]  = eta_sum_out_tmp[1][18];
        eta_sum[1][4]  = eta_sum_out_tmp[1][19];
        eta_sum[1][5]  = eta_sum_out_tmp[1][20];
        eta_sum[1][6]  = eta_sum_out_tmp[1][21];
        eta_sum[1][7]  = eta_sum_out_tmp[1][22];
        eta_sum[1][8]  = eta_sum_out_tmp[1][23];
        eta_sum[1][9]  = eta_sum_out_tmp[1][24];
        eta_sum[1][10]  = eta_sum_out_tmp[1][25];
        eta_sum[1][11]  = eta_sum_out_tmp[1][26];
        eta_sum[1][12]  = eta_sum_out_tmp[1][27];
        eta_sum[1][13]  = eta_sum_out_tmp[1][28];
        eta_sum[1][14]  = eta_sum_out_tmp[1][29];
        eta_sum[1][15]  = eta_sum_out_tmp[1][30];
        eta_sum[1][16]  = eta_sum_out_tmp[1][31];
        eta_sum[1][17]  = eta_sum_out_tmp[1][32];
        eta_sum[1][18]  = eta_sum_out_tmp[1][33];
        eta_sum[1][19]  = eta_sum_out_tmp[1][34];
        eta_sum[1][20]  = eta_sum_out_tmp[1][35];
        eta_sum[1][21]  = eta_sum_out_tmp[1][36];
        eta_sum[1][22]  = eta_sum_out_tmp[1][37];
        eta_sum[1][23]  = eta_sum_out_tmp[1][38];
        eta_sum[1][24]  = eta_sum_out_tmp[1][39];
        eta_sum[1][25]  = eta_sum_out_tmp[1][40];
        eta_sum[1][26]  = eta_sum_out_tmp[1][41];
    end
 
    4:begin 
        eta_sum[1][0]  = eta_sum_out_tmp[1][0];
        eta_sum[1][1]  = eta_sum_out_tmp[1][1];
        eta_sum[1][2]  = eta_sum_out_tmp[1][2];
        eta_sum[1][3]  = eta_sum_out_tmp[1][3];
        eta_sum[1][4]  = eta_sum_out_tmp[1][4];
        eta_sum[1][5]  = eta_sum_out_tmp[1][5];
        eta_sum[1][6]  = eta_sum_out_tmp[1][6];
        eta_sum[1][7]  = eta_sum_out_tmp[1][7];
        eta_sum[1][8]  = eta_sum_out_tmp[1][8];
        eta_sum[1][9]  = eta_sum_out_tmp[1][9];
        eta_sum[1][10]  = eta_sum_out_tmp[1][10];
        eta_sum[1][11]  = eta_sum_out_tmp[1][11];
        eta_sum[1][12]  = eta_sum_out_tmp[1][12];
        eta_sum[1][13]  = eta_sum_out_tmp[1][13];
        eta_sum[1][14]  = eta_sum_out_tmp[1][14];
        eta_sum[1][15]  = eta_sum_out_tmp[1][15];
        eta_sum[1][16]  = eta_sum_out_tmp[1][16];
        eta_sum[1][17]  = eta_sum_out_tmp[1][17];
        eta_sum[1][18]  = eta_sum_out_tmp[1][18];
        eta_sum[1][19]  = eta_sum_out_tmp[1][19];
        eta_sum[1][20]  = eta_sum_out_tmp[1][20];
        eta_sum[1][21]  = eta_sum_out_tmp[1][21];
        eta_sum[1][22]  = eta_sum_out_tmp[1][22];
        eta_sum[1][23]  = eta_sum_out_tmp[1][23];
        eta_sum[1][24]  = eta_sum_out_tmp[1][24];
        eta_sum[1][25]  = eta_sum_out_tmp[1][25];
        eta_sum[1][26]  = eta_sum_out_tmp[1][26];
        eta_sum[1][27]  = eta_sum_out_tmp[1][27];
        eta_sum[1][28]  = eta_sum_out_tmp[1][28];
        eta_sum[1][29]  = eta_sum_out_tmp[1][29];
        eta_sum[1][30]  = eta_sum_out_tmp[1][30];
        eta_sum[1][31]  = eta_sum_out_tmp[1][31];
        eta_sum[1][32]  = eta_sum_out_tmp[1][32];
        eta_sum[1][33]  = eta_sum_out_tmp[1][33];
        eta_sum[1][34]  = eta_sum_out_tmp[1][34];
        eta_sum[1][35]  = eta_sum_out_tmp[1][35];
        eta_sum[1][36]  = eta_sum_out_tmp[1][36];
        eta_sum[1][37]  = eta_sum_out_tmp[1][37];
        eta_sum[1][38]  = eta_sum_out_tmp[1][38];
        eta_sum[1][39]  = eta_sum_out_tmp[1][39];
        eta_sum[1][40]  = eta_sum_out_tmp[1][40];
        eta_sum[1][41]  = eta_sum_out_tmp[1][41];
    end
 
    5:begin 
        eta_sum[1][0]  = eta_sum_out_tmp[1][0];
        eta_sum[1][1]  = eta_sum_out_tmp[1][1];
        eta_sum[1][2]  = eta_sum_out_tmp[1][2];
        eta_sum[1][3]  = eta_sum_out_tmp[1][3];
        eta_sum[1][4]  = eta_sum_out_tmp[1][4];
        eta_sum[1][5]  = eta_sum_out_tmp[1][5];
        eta_sum[1][6]  = eta_sum_out_tmp[1][6];
        eta_sum[1][7]  = eta_sum_out_tmp[1][7];
        eta_sum[1][8]  = eta_sum_out_tmp[1][8];
        eta_sum[1][9]  = eta_sum_out_tmp[1][9];
        eta_sum[1][10]  = eta_sum_out_tmp[1][10];
        eta_sum[1][11]  = eta_sum_out_tmp[1][11];
        eta_sum[1][12]  = eta_sum_out_tmp[1][12];
        eta_sum[1][13]  = eta_sum_out_tmp[1][13];
        eta_sum[1][14]  = eta_sum_out_tmp[1][14];
        eta_sum[1][15]  = eta_sum_out_tmp[1][15];
        eta_sum[1][16]  = eta_sum_out_tmp[1][16];
        eta_sum[1][17]  = eta_sum_out_tmp[1][17];
        eta_sum[1][18]  = eta_sum_out_tmp[1][18];
        eta_sum[1][19]  = eta_sum_out_tmp[1][19];
        eta_sum[1][20]  = eta_sum_out_tmp[1][20];
        eta_sum[1][21]  = eta_sum_out_tmp[1][21];
        eta_sum[1][22]  = eta_sum_out_tmp[1][22];
        eta_sum[1][23]  = eta_sum_out_tmp[1][23];
        eta_sum[1][24]  = eta_sum_out_tmp[1][24];
        eta_sum[1][25]  = eta_sum_out_tmp[1][25];
        eta_sum[1][26]  = eta_sum_out_tmp[1][26];
        eta_sum[1][27]  = eta_sum_out_tmp[1][27];
        eta_sum[1][28]  = eta_sum_out_tmp[1][28];
        eta_sum[1][29]  = eta_sum_out_tmp[1][29];
        eta_sum[1][30]  = eta_sum_out_tmp[1][30];
        eta_sum[1][31]  = eta_sum_out_tmp[1][31];
        eta_sum[1][32]  = eta_sum_out_tmp[1][32];
        eta_sum[1][33]  = eta_sum_out_tmp[1][33];
        eta_sum[1][34]  = eta_sum_out_tmp[1][34];
        eta_sum[1][35]  = eta_sum_out_tmp[1][35];
        eta_sum[1][36]  = eta_sum_out_tmp[1][36];
        eta_sum[1][37]  = eta_sum_out_tmp[1][37];
        eta_sum[1][38]  = eta_sum_out_tmp[1][38];
        eta_sum[1][39]  = eta_sum_out_tmp[1][39];
        eta_sum[1][40]  = eta_sum_out_tmp[1][40];
        eta_sum[1][41]  = eta_sum_out_tmp[1][41];
    end
 
    6:begin 
        eta_sum[1][31]  = eta_sum_out_tmp[1][0];
        eta_sum[1][32]  = eta_sum_out_tmp[1][1];
        eta_sum[1][33]  = eta_sum_out_tmp[1][2];
        eta_sum[1][34]  = eta_sum_out_tmp[1][3];
        eta_sum[1][35]  = eta_sum_out_tmp[1][4];
        eta_sum[1][36]  = eta_sum_out_tmp[1][5];
        eta_sum[1][37]  = eta_sum_out_tmp[1][6];
        eta_sum[1][38]  = eta_sum_out_tmp[1][7];
        eta_sum[1][39]  = eta_sum_out_tmp[1][8];
        eta_sum[1][40]  = eta_sum_out_tmp[1][9];
        eta_sum[1][41]  = eta_sum_out_tmp[1][10];
        eta_sum[1][0]  = eta_sum_out_tmp[1][11];
        eta_sum[1][1]  = eta_sum_out_tmp[1][12];
        eta_sum[1][2]  = eta_sum_out_tmp[1][13];
        eta_sum[1][3]  = eta_sum_out_tmp[1][14];
        eta_sum[1][4]  = eta_sum_out_tmp[1][15];
        eta_sum[1][5]  = eta_sum_out_tmp[1][16];
        eta_sum[1][6]  = eta_sum_out_tmp[1][17];
        eta_sum[1][7]  = eta_sum_out_tmp[1][18];
        eta_sum[1][8]  = eta_sum_out_tmp[1][19];
        eta_sum[1][9]  = eta_sum_out_tmp[1][20];
        eta_sum[1][10]  = eta_sum_out_tmp[1][21];
        eta_sum[1][11]  = eta_sum_out_tmp[1][22];
        eta_sum[1][12]  = eta_sum_out_tmp[1][23];
        eta_sum[1][13]  = eta_sum_out_tmp[1][24];
        eta_sum[1][14]  = eta_sum_out_tmp[1][25];
        eta_sum[1][15]  = eta_sum_out_tmp[1][26];
        eta_sum[1][16]  = eta_sum_out_tmp[1][27];
        eta_sum[1][17]  = eta_sum_out_tmp[1][28];
        eta_sum[1][18]  = eta_sum_out_tmp[1][29];
        eta_sum[1][19]  = eta_sum_out_tmp[1][30];
        eta_sum[1][20]  = eta_sum_out_tmp[1][31];
        eta_sum[1][21]  = eta_sum_out_tmp[1][32];
        eta_sum[1][22]  = eta_sum_out_tmp[1][33];
        eta_sum[1][23]  = eta_sum_out_tmp[1][34];
        eta_sum[1][24]  = eta_sum_out_tmp[1][35];
        eta_sum[1][25]  = eta_sum_out_tmp[1][36];
        eta_sum[1][26]  = eta_sum_out_tmp[1][37];
        eta_sum[1][27]  = eta_sum_out_tmp[1][38];
        eta_sum[1][28]  = eta_sum_out_tmp[1][39];
        eta_sum[1][29]  = eta_sum_out_tmp[1][40];
        eta_sum[1][30]  = eta_sum_out_tmp[1][41];
    end
 
    7:begin 
        eta_sum[1][22]  = eta_sum_out_tmp[1][0];
        eta_sum[1][23]  = eta_sum_out_tmp[1][1];
        eta_sum[1][24]  = eta_sum_out_tmp[1][2];
        eta_sum[1][25]  = eta_sum_out_tmp[1][3];
        eta_sum[1][26]  = eta_sum_out_tmp[1][4];
        eta_sum[1][27]  = eta_sum_out_tmp[1][5];
        eta_sum[1][28]  = eta_sum_out_tmp[1][6];
        eta_sum[1][29]  = eta_sum_out_tmp[1][7];
        eta_sum[1][30]  = eta_sum_out_tmp[1][8];
        eta_sum[1][31]  = eta_sum_out_tmp[1][9];
        eta_sum[1][32]  = eta_sum_out_tmp[1][10];
        eta_sum[1][33]  = eta_sum_out_tmp[1][11];
        eta_sum[1][34]  = eta_sum_out_tmp[1][12];
        eta_sum[1][35]  = eta_sum_out_tmp[1][13];
        eta_sum[1][36]  = eta_sum_out_tmp[1][14];
        eta_sum[1][37]  = eta_sum_out_tmp[1][15];
        eta_sum[1][38]  = eta_sum_out_tmp[1][16];
        eta_sum[1][39]  = eta_sum_out_tmp[1][17];
        eta_sum[1][40]  = eta_sum_out_tmp[1][18];
        eta_sum[1][41]  = eta_sum_out_tmp[1][19];
        eta_sum[1][0]  = eta_sum_out_tmp[1][20];
        eta_sum[1][1]  = eta_sum_out_tmp[1][21];
        eta_sum[1][2]  = eta_sum_out_tmp[1][22];
        eta_sum[1][3]  = eta_sum_out_tmp[1][23];
        eta_sum[1][4]  = eta_sum_out_tmp[1][24];
        eta_sum[1][5]  = eta_sum_out_tmp[1][25];
        eta_sum[1][6]  = eta_sum_out_tmp[1][26];
        eta_sum[1][7]  = eta_sum_out_tmp[1][27];
        eta_sum[1][8]  = eta_sum_out_tmp[1][28];
        eta_sum[1][9]  = eta_sum_out_tmp[1][29];
        eta_sum[1][10]  = eta_sum_out_tmp[1][30];
        eta_sum[1][11]  = eta_sum_out_tmp[1][31];
        eta_sum[1][12]  = eta_sum_out_tmp[1][32];
        eta_sum[1][13]  = eta_sum_out_tmp[1][33];
        eta_sum[1][14]  = eta_sum_out_tmp[1][34];
        eta_sum[1][15]  = eta_sum_out_tmp[1][35];
        eta_sum[1][16]  = eta_sum_out_tmp[1][36];
        eta_sum[1][17]  = eta_sum_out_tmp[1][37];
        eta_sum[1][18]  = eta_sum_out_tmp[1][38];
        eta_sum[1][19]  = eta_sum_out_tmp[1][39];
        eta_sum[1][20]  = eta_sum_out_tmp[1][40];
        eta_sum[1][21]  = eta_sum_out_tmp[1][41];
    end
 
endcase
end

if (chk_n_output_valid[0] & active_cols[2]) begin
case (curr_layer)
    0:begin 
        eta_sum[2][38]  = eta_sum_out_tmp[2][0];
        eta_sum[2][39]  = eta_sum_out_tmp[2][1];
        eta_sum[2][40]  = eta_sum_out_tmp[2][2];
        eta_sum[2][41]  = eta_sum_out_tmp[2][3];
        eta_sum[2][0]  = eta_sum_out_tmp[2][4];
        eta_sum[2][1]  = eta_sum_out_tmp[2][5];
        eta_sum[2][2]  = eta_sum_out_tmp[2][6];
        eta_sum[2][3]  = eta_sum_out_tmp[2][7];
        eta_sum[2][4]  = eta_sum_out_tmp[2][8];
        eta_sum[2][5]  = eta_sum_out_tmp[2][9];
        eta_sum[2][6]  = eta_sum_out_tmp[2][10];
        eta_sum[2][7]  = eta_sum_out_tmp[2][11];
        eta_sum[2][8]  = eta_sum_out_tmp[2][12];
        eta_sum[2][9]  = eta_sum_out_tmp[2][13];
        eta_sum[2][10]  = eta_sum_out_tmp[2][14];
        eta_sum[2][11]  = eta_sum_out_tmp[2][15];
        eta_sum[2][12]  = eta_sum_out_tmp[2][16];
        eta_sum[2][13]  = eta_sum_out_tmp[2][17];
        eta_sum[2][14]  = eta_sum_out_tmp[2][18];
        eta_sum[2][15]  = eta_sum_out_tmp[2][19];
        eta_sum[2][16]  = eta_sum_out_tmp[2][20];
        eta_sum[2][17]  = eta_sum_out_tmp[2][21];
        eta_sum[2][18]  = eta_sum_out_tmp[2][22];
        eta_sum[2][19]  = eta_sum_out_tmp[2][23];
        eta_sum[2][20]  = eta_sum_out_tmp[2][24];
        eta_sum[2][21]  = eta_sum_out_tmp[2][25];
        eta_sum[2][22]  = eta_sum_out_tmp[2][26];
        eta_sum[2][23]  = eta_sum_out_tmp[2][27];
        eta_sum[2][24]  = eta_sum_out_tmp[2][28];
        eta_sum[2][25]  = eta_sum_out_tmp[2][29];
        eta_sum[2][26]  = eta_sum_out_tmp[2][30];
        eta_sum[2][27]  = eta_sum_out_tmp[2][31];
        eta_sum[2][28]  = eta_sum_out_tmp[2][32];
        eta_sum[2][29]  = eta_sum_out_tmp[2][33];
        eta_sum[2][30]  = eta_sum_out_tmp[2][34];
        eta_sum[2][31]  = eta_sum_out_tmp[2][35];
        eta_sum[2][32]  = eta_sum_out_tmp[2][36];
        eta_sum[2][33]  = eta_sum_out_tmp[2][37];
        eta_sum[2][34]  = eta_sum_out_tmp[2][38];
        eta_sum[2][35]  = eta_sum_out_tmp[2][39];
        eta_sum[2][36]  = eta_sum_out_tmp[2][40];
        eta_sum[2][37]  = eta_sum_out_tmp[2][41];
    end
 
    1:begin 
        eta_sum[2][35]  = eta_sum_out_tmp[2][0];
        eta_sum[2][36]  = eta_sum_out_tmp[2][1];
        eta_sum[2][37]  = eta_sum_out_tmp[2][2];
        eta_sum[2][38]  = eta_sum_out_tmp[2][3];
        eta_sum[2][39]  = eta_sum_out_tmp[2][4];
        eta_sum[2][40]  = eta_sum_out_tmp[2][5];
        eta_sum[2][41]  = eta_sum_out_tmp[2][6];
        eta_sum[2][0]  = eta_sum_out_tmp[2][7];
        eta_sum[2][1]  = eta_sum_out_tmp[2][8];
        eta_sum[2][2]  = eta_sum_out_tmp[2][9];
        eta_sum[2][3]  = eta_sum_out_tmp[2][10];
        eta_sum[2][4]  = eta_sum_out_tmp[2][11];
        eta_sum[2][5]  = eta_sum_out_tmp[2][12];
        eta_sum[2][6]  = eta_sum_out_tmp[2][13];
        eta_sum[2][7]  = eta_sum_out_tmp[2][14];
        eta_sum[2][8]  = eta_sum_out_tmp[2][15];
        eta_sum[2][9]  = eta_sum_out_tmp[2][16];
        eta_sum[2][10]  = eta_sum_out_tmp[2][17];
        eta_sum[2][11]  = eta_sum_out_tmp[2][18];
        eta_sum[2][12]  = eta_sum_out_tmp[2][19];
        eta_sum[2][13]  = eta_sum_out_tmp[2][20];
        eta_sum[2][14]  = eta_sum_out_tmp[2][21];
        eta_sum[2][15]  = eta_sum_out_tmp[2][22];
        eta_sum[2][16]  = eta_sum_out_tmp[2][23];
        eta_sum[2][17]  = eta_sum_out_tmp[2][24];
        eta_sum[2][18]  = eta_sum_out_tmp[2][25];
        eta_sum[2][19]  = eta_sum_out_tmp[2][26];
        eta_sum[2][20]  = eta_sum_out_tmp[2][27];
        eta_sum[2][21]  = eta_sum_out_tmp[2][28];
        eta_sum[2][22]  = eta_sum_out_tmp[2][29];
        eta_sum[2][23]  = eta_sum_out_tmp[2][30];
        eta_sum[2][24]  = eta_sum_out_tmp[2][31];
        eta_sum[2][25]  = eta_sum_out_tmp[2][32];
        eta_sum[2][26]  = eta_sum_out_tmp[2][33];
        eta_sum[2][27]  = eta_sum_out_tmp[2][34];
        eta_sum[2][28]  = eta_sum_out_tmp[2][35];
        eta_sum[2][29]  = eta_sum_out_tmp[2][36];
        eta_sum[2][30]  = eta_sum_out_tmp[2][37];
        eta_sum[2][31]  = eta_sum_out_tmp[2][38];
        eta_sum[2][32]  = eta_sum_out_tmp[2][39];
        eta_sum[2][33]  = eta_sum_out_tmp[2][40];
        eta_sum[2][34]  = eta_sum_out_tmp[2][41];
    end
 
    2:begin 
        eta_sum[2][0]  = eta_sum_out_tmp[2][0];
        eta_sum[2][1]  = eta_sum_out_tmp[2][1];
        eta_sum[2][2]  = eta_sum_out_tmp[2][2];
        eta_sum[2][3]  = eta_sum_out_tmp[2][3];
        eta_sum[2][4]  = eta_sum_out_tmp[2][4];
        eta_sum[2][5]  = eta_sum_out_tmp[2][5];
        eta_sum[2][6]  = eta_sum_out_tmp[2][6];
        eta_sum[2][7]  = eta_sum_out_tmp[2][7];
        eta_sum[2][8]  = eta_sum_out_tmp[2][8];
        eta_sum[2][9]  = eta_sum_out_tmp[2][9];
        eta_sum[2][10]  = eta_sum_out_tmp[2][10];
        eta_sum[2][11]  = eta_sum_out_tmp[2][11];
        eta_sum[2][12]  = eta_sum_out_tmp[2][12];
        eta_sum[2][13]  = eta_sum_out_tmp[2][13];
        eta_sum[2][14]  = eta_sum_out_tmp[2][14];
        eta_sum[2][15]  = eta_sum_out_tmp[2][15];
        eta_sum[2][16]  = eta_sum_out_tmp[2][16];
        eta_sum[2][17]  = eta_sum_out_tmp[2][17];
        eta_sum[2][18]  = eta_sum_out_tmp[2][18];
        eta_sum[2][19]  = eta_sum_out_tmp[2][19];
        eta_sum[2][20]  = eta_sum_out_tmp[2][20];
        eta_sum[2][21]  = eta_sum_out_tmp[2][21];
        eta_sum[2][22]  = eta_sum_out_tmp[2][22];
        eta_sum[2][23]  = eta_sum_out_tmp[2][23];
        eta_sum[2][24]  = eta_sum_out_tmp[2][24];
        eta_sum[2][25]  = eta_sum_out_tmp[2][25];
        eta_sum[2][26]  = eta_sum_out_tmp[2][26];
        eta_sum[2][27]  = eta_sum_out_tmp[2][27];
        eta_sum[2][28]  = eta_sum_out_tmp[2][28];
        eta_sum[2][29]  = eta_sum_out_tmp[2][29];
        eta_sum[2][30]  = eta_sum_out_tmp[2][30];
        eta_sum[2][31]  = eta_sum_out_tmp[2][31];
        eta_sum[2][32]  = eta_sum_out_tmp[2][32];
        eta_sum[2][33]  = eta_sum_out_tmp[2][33];
        eta_sum[2][34]  = eta_sum_out_tmp[2][34];
        eta_sum[2][35]  = eta_sum_out_tmp[2][35];
        eta_sum[2][36]  = eta_sum_out_tmp[2][36];
        eta_sum[2][37]  = eta_sum_out_tmp[2][37];
        eta_sum[2][38]  = eta_sum_out_tmp[2][38];
        eta_sum[2][39]  = eta_sum_out_tmp[2][39];
        eta_sum[2][40]  = eta_sum_out_tmp[2][40];
        eta_sum[2][41]  = eta_sum_out_tmp[2][41];
    end
 
    3:begin 
        eta_sum[2][0]  = eta_sum_out_tmp[2][0];
        eta_sum[2][1]  = eta_sum_out_tmp[2][1];
        eta_sum[2][2]  = eta_sum_out_tmp[2][2];
        eta_sum[2][3]  = eta_sum_out_tmp[2][3];
        eta_sum[2][4]  = eta_sum_out_tmp[2][4];
        eta_sum[2][5]  = eta_sum_out_tmp[2][5];
        eta_sum[2][6]  = eta_sum_out_tmp[2][6];
        eta_sum[2][7]  = eta_sum_out_tmp[2][7];
        eta_sum[2][8]  = eta_sum_out_tmp[2][8];
        eta_sum[2][9]  = eta_sum_out_tmp[2][9];
        eta_sum[2][10]  = eta_sum_out_tmp[2][10];
        eta_sum[2][11]  = eta_sum_out_tmp[2][11];
        eta_sum[2][12]  = eta_sum_out_tmp[2][12];
        eta_sum[2][13]  = eta_sum_out_tmp[2][13];
        eta_sum[2][14]  = eta_sum_out_tmp[2][14];
        eta_sum[2][15]  = eta_sum_out_tmp[2][15];
        eta_sum[2][16]  = eta_sum_out_tmp[2][16];
        eta_sum[2][17]  = eta_sum_out_tmp[2][17];
        eta_sum[2][18]  = eta_sum_out_tmp[2][18];
        eta_sum[2][19]  = eta_sum_out_tmp[2][19];
        eta_sum[2][20]  = eta_sum_out_tmp[2][20];
        eta_sum[2][21]  = eta_sum_out_tmp[2][21];
        eta_sum[2][22]  = eta_sum_out_tmp[2][22];
        eta_sum[2][23]  = eta_sum_out_tmp[2][23];
        eta_sum[2][24]  = eta_sum_out_tmp[2][24];
        eta_sum[2][25]  = eta_sum_out_tmp[2][25];
        eta_sum[2][26]  = eta_sum_out_tmp[2][26];
        eta_sum[2][27]  = eta_sum_out_tmp[2][27];
        eta_sum[2][28]  = eta_sum_out_tmp[2][28];
        eta_sum[2][29]  = eta_sum_out_tmp[2][29];
        eta_sum[2][30]  = eta_sum_out_tmp[2][30];
        eta_sum[2][31]  = eta_sum_out_tmp[2][31];
        eta_sum[2][32]  = eta_sum_out_tmp[2][32];
        eta_sum[2][33]  = eta_sum_out_tmp[2][33];
        eta_sum[2][34]  = eta_sum_out_tmp[2][34];
        eta_sum[2][35]  = eta_sum_out_tmp[2][35];
        eta_sum[2][36]  = eta_sum_out_tmp[2][36];
        eta_sum[2][37]  = eta_sum_out_tmp[2][37];
        eta_sum[2][38]  = eta_sum_out_tmp[2][38];
        eta_sum[2][39]  = eta_sum_out_tmp[2][39];
        eta_sum[2][40]  = eta_sum_out_tmp[2][40];
        eta_sum[2][41]  = eta_sum_out_tmp[2][41];
    end
 
    4:begin 
        eta_sum[2][41]  = eta_sum_out_tmp[2][0];
        eta_sum[2][0]  = eta_sum_out_tmp[2][1];
        eta_sum[2][1]  = eta_sum_out_tmp[2][2];
        eta_sum[2][2]  = eta_sum_out_tmp[2][3];
        eta_sum[2][3]  = eta_sum_out_tmp[2][4];
        eta_sum[2][4]  = eta_sum_out_tmp[2][5];
        eta_sum[2][5]  = eta_sum_out_tmp[2][6];
        eta_sum[2][6]  = eta_sum_out_tmp[2][7];
        eta_sum[2][7]  = eta_sum_out_tmp[2][8];
        eta_sum[2][8]  = eta_sum_out_tmp[2][9];
        eta_sum[2][9]  = eta_sum_out_tmp[2][10];
        eta_sum[2][10]  = eta_sum_out_tmp[2][11];
        eta_sum[2][11]  = eta_sum_out_tmp[2][12];
        eta_sum[2][12]  = eta_sum_out_tmp[2][13];
        eta_sum[2][13]  = eta_sum_out_tmp[2][14];
        eta_sum[2][14]  = eta_sum_out_tmp[2][15];
        eta_sum[2][15]  = eta_sum_out_tmp[2][16];
        eta_sum[2][16]  = eta_sum_out_tmp[2][17];
        eta_sum[2][17]  = eta_sum_out_tmp[2][18];
        eta_sum[2][18]  = eta_sum_out_tmp[2][19];
        eta_sum[2][19]  = eta_sum_out_tmp[2][20];
        eta_sum[2][20]  = eta_sum_out_tmp[2][21];
        eta_sum[2][21]  = eta_sum_out_tmp[2][22];
        eta_sum[2][22]  = eta_sum_out_tmp[2][23];
        eta_sum[2][23]  = eta_sum_out_tmp[2][24];
        eta_sum[2][24]  = eta_sum_out_tmp[2][25];
        eta_sum[2][25]  = eta_sum_out_tmp[2][26];
        eta_sum[2][26]  = eta_sum_out_tmp[2][27];
        eta_sum[2][27]  = eta_sum_out_tmp[2][28];
        eta_sum[2][28]  = eta_sum_out_tmp[2][29];
        eta_sum[2][29]  = eta_sum_out_tmp[2][30];
        eta_sum[2][30]  = eta_sum_out_tmp[2][31];
        eta_sum[2][31]  = eta_sum_out_tmp[2][32];
        eta_sum[2][32]  = eta_sum_out_tmp[2][33];
        eta_sum[2][33]  = eta_sum_out_tmp[2][34];
        eta_sum[2][34]  = eta_sum_out_tmp[2][35];
        eta_sum[2][35]  = eta_sum_out_tmp[2][36];
        eta_sum[2][36]  = eta_sum_out_tmp[2][37];
        eta_sum[2][37]  = eta_sum_out_tmp[2][38];
        eta_sum[2][38]  = eta_sum_out_tmp[2][39];
        eta_sum[2][39]  = eta_sum_out_tmp[2][40];
        eta_sum[2][40]  = eta_sum_out_tmp[2][41];
    end
 
    5:begin 
        eta_sum[2][0]  = eta_sum_out_tmp[2][0];
        eta_sum[2][1]  = eta_sum_out_tmp[2][1];
        eta_sum[2][2]  = eta_sum_out_tmp[2][2];
        eta_sum[2][3]  = eta_sum_out_tmp[2][3];
        eta_sum[2][4]  = eta_sum_out_tmp[2][4];
        eta_sum[2][5]  = eta_sum_out_tmp[2][5];
        eta_sum[2][6]  = eta_sum_out_tmp[2][6];
        eta_sum[2][7]  = eta_sum_out_tmp[2][7];
        eta_sum[2][8]  = eta_sum_out_tmp[2][8];
        eta_sum[2][9]  = eta_sum_out_tmp[2][9];
        eta_sum[2][10]  = eta_sum_out_tmp[2][10];
        eta_sum[2][11]  = eta_sum_out_tmp[2][11];
        eta_sum[2][12]  = eta_sum_out_tmp[2][12];
        eta_sum[2][13]  = eta_sum_out_tmp[2][13];
        eta_sum[2][14]  = eta_sum_out_tmp[2][14];
        eta_sum[2][15]  = eta_sum_out_tmp[2][15];
        eta_sum[2][16]  = eta_sum_out_tmp[2][16];
        eta_sum[2][17]  = eta_sum_out_tmp[2][17];
        eta_sum[2][18]  = eta_sum_out_tmp[2][18];
        eta_sum[2][19]  = eta_sum_out_tmp[2][19];
        eta_sum[2][20]  = eta_sum_out_tmp[2][20];
        eta_sum[2][21]  = eta_sum_out_tmp[2][21];
        eta_sum[2][22]  = eta_sum_out_tmp[2][22];
        eta_sum[2][23]  = eta_sum_out_tmp[2][23];
        eta_sum[2][24]  = eta_sum_out_tmp[2][24];
        eta_sum[2][25]  = eta_sum_out_tmp[2][25];
        eta_sum[2][26]  = eta_sum_out_tmp[2][26];
        eta_sum[2][27]  = eta_sum_out_tmp[2][27];
        eta_sum[2][28]  = eta_sum_out_tmp[2][28];
        eta_sum[2][29]  = eta_sum_out_tmp[2][29];
        eta_sum[2][30]  = eta_sum_out_tmp[2][30];
        eta_sum[2][31]  = eta_sum_out_tmp[2][31];
        eta_sum[2][32]  = eta_sum_out_tmp[2][32];
        eta_sum[2][33]  = eta_sum_out_tmp[2][33];
        eta_sum[2][34]  = eta_sum_out_tmp[2][34];
        eta_sum[2][35]  = eta_sum_out_tmp[2][35];
        eta_sum[2][36]  = eta_sum_out_tmp[2][36];
        eta_sum[2][37]  = eta_sum_out_tmp[2][37];
        eta_sum[2][38]  = eta_sum_out_tmp[2][38];
        eta_sum[2][39]  = eta_sum_out_tmp[2][39];
        eta_sum[2][40]  = eta_sum_out_tmp[2][40];
        eta_sum[2][41]  = eta_sum_out_tmp[2][41];
    end
 
    6:begin 
        eta_sum[2][0]  = eta_sum_out_tmp[2][0];
        eta_sum[2][1]  = eta_sum_out_tmp[2][1];
        eta_sum[2][2]  = eta_sum_out_tmp[2][2];
        eta_sum[2][3]  = eta_sum_out_tmp[2][3];
        eta_sum[2][4]  = eta_sum_out_tmp[2][4];
        eta_sum[2][5]  = eta_sum_out_tmp[2][5];
        eta_sum[2][6]  = eta_sum_out_tmp[2][6];
        eta_sum[2][7]  = eta_sum_out_tmp[2][7];
        eta_sum[2][8]  = eta_sum_out_tmp[2][8];
        eta_sum[2][9]  = eta_sum_out_tmp[2][9];
        eta_sum[2][10]  = eta_sum_out_tmp[2][10];
        eta_sum[2][11]  = eta_sum_out_tmp[2][11];
        eta_sum[2][12]  = eta_sum_out_tmp[2][12];
        eta_sum[2][13]  = eta_sum_out_tmp[2][13];
        eta_sum[2][14]  = eta_sum_out_tmp[2][14];
        eta_sum[2][15]  = eta_sum_out_tmp[2][15];
        eta_sum[2][16]  = eta_sum_out_tmp[2][16];
        eta_sum[2][17]  = eta_sum_out_tmp[2][17];
        eta_sum[2][18]  = eta_sum_out_tmp[2][18];
        eta_sum[2][19]  = eta_sum_out_tmp[2][19];
        eta_sum[2][20]  = eta_sum_out_tmp[2][20];
        eta_sum[2][21]  = eta_sum_out_tmp[2][21];
        eta_sum[2][22]  = eta_sum_out_tmp[2][22];
        eta_sum[2][23]  = eta_sum_out_tmp[2][23];
        eta_sum[2][24]  = eta_sum_out_tmp[2][24];
        eta_sum[2][25]  = eta_sum_out_tmp[2][25];
        eta_sum[2][26]  = eta_sum_out_tmp[2][26];
        eta_sum[2][27]  = eta_sum_out_tmp[2][27];
        eta_sum[2][28]  = eta_sum_out_tmp[2][28];
        eta_sum[2][29]  = eta_sum_out_tmp[2][29];
        eta_sum[2][30]  = eta_sum_out_tmp[2][30];
        eta_sum[2][31]  = eta_sum_out_tmp[2][31];
        eta_sum[2][32]  = eta_sum_out_tmp[2][32];
        eta_sum[2][33]  = eta_sum_out_tmp[2][33];
        eta_sum[2][34]  = eta_sum_out_tmp[2][34];
        eta_sum[2][35]  = eta_sum_out_tmp[2][35];
        eta_sum[2][36]  = eta_sum_out_tmp[2][36];
        eta_sum[2][37]  = eta_sum_out_tmp[2][37];
        eta_sum[2][38]  = eta_sum_out_tmp[2][38];
        eta_sum[2][39]  = eta_sum_out_tmp[2][39];
        eta_sum[2][40]  = eta_sum_out_tmp[2][40];
        eta_sum[2][41]  = eta_sum_out_tmp[2][41];
    end
 
    7:begin 
        eta_sum[2][0]  = eta_sum_out_tmp[2][0];
        eta_sum[2][1]  = eta_sum_out_tmp[2][1];
        eta_sum[2][2]  = eta_sum_out_tmp[2][2];
        eta_sum[2][3]  = eta_sum_out_tmp[2][3];
        eta_sum[2][4]  = eta_sum_out_tmp[2][4];
        eta_sum[2][5]  = eta_sum_out_tmp[2][5];
        eta_sum[2][6]  = eta_sum_out_tmp[2][6];
        eta_sum[2][7]  = eta_sum_out_tmp[2][7];
        eta_sum[2][8]  = eta_sum_out_tmp[2][8];
        eta_sum[2][9]  = eta_sum_out_tmp[2][9];
        eta_sum[2][10]  = eta_sum_out_tmp[2][10];
        eta_sum[2][11]  = eta_sum_out_tmp[2][11];
        eta_sum[2][12]  = eta_sum_out_tmp[2][12];
        eta_sum[2][13]  = eta_sum_out_tmp[2][13];
        eta_sum[2][14]  = eta_sum_out_tmp[2][14];
        eta_sum[2][15]  = eta_sum_out_tmp[2][15];
        eta_sum[2][16]  = eta_sum_out_tmp[2][16];
        eta_sum[2][17]  = eta_sum_out_tmp[2][17];
        eta_sum[2][18]  = eta_sum_out_tmp[2][18];
        eta_sum[2][19]  = eta_sum_out_tmp[2][19];
        eta_sum[2][20]  = eta_sum_out_tmp[2][20];
        eta_sum[2][21]  = eta_sum_out_tmp[2][21];
        eta_sum[2][22]  = eta_sum_out_tmp[2][22];
        eta_sum[2][23]  = eta_sum_out_tmp[2][23];
        eta_sum[2][24]  = eta_sum_out_tmp[2][24];
        eta_sum[2][25]  = eta_sum_out_tmp[2][25];
        eta_sum[2][26]  = eta_sum_out_tmp[2][26];
        eta_sum[2][27]  = eta_sum_out_tmp[2][27];
        eta_sum[2][28]  = eta_sum_out_tmp[2][28];
        eta_sum[2][29]  = eta_sum_out_tmp[2][29];
        eta_sum[2][30]  = eta_sum_out_tmp[2][30];
        eta_sum[2][31]  = eta_sum_out_tmp[2][31];
        eta_sum[2][32]  = eta_sum_out_tmp[2][32];
        eta_sum[2][33]  = eta_sum_out_tmp[2][33];
        eta_sum[2][34]  = eta_sum_out_tmp[2][34];
        eta_sum[2][35]  = eta_sum_out_tmp[2][35];
        eta_sum[2][36]  = eta_sum_out_tmp[2][36];
        eta_sum[2][37]  = eta_sum_out_tmp[2][37];
        eta_sum[2][38]  = eta_sum_out_tmp[2][38];
        eta_sum[2][39]  = eta_sum_out_tmp[2][39];
        eta_sum[2][40]  = eta_sum_out_tmp[2][40];
        eta_sum[2][41]  = eta_sum_out_tmp[2][41];
    end
 
endcase
end

if (chk_n_output_valid[0] & active_cols[3]) begin
case (curr_layer)
    0:begin 
        eta_sum[3][0]  = eta_sum_out_tmp[3][0];
        eta_sum[3][1]  = eta_sum_out_tmp[3][1];
        eta_sum[3][2]  = eta_sum_out_tmp[3][2];
        eta_sum[3][3]  = eta_sum_out_tmp[3][3];
        eta_sum[3][4]  = eta_sum_out_tmp[3][4];
        eta_sum[3][5]  = eta_sum_out_tmp[3][5];
        eta_sum[3][6]  = eta_sum_out_tmp[3][6];
        eta_sum[3][7]  = eta_sum_out_tmp[3][7];
        eta_sum[3][8]  = eta_sum_out_tmp[3][8];
        eta_sum[3][9]  = eta_sum_out_tmp[3][9];
        eta_sum[3][10]  = eta_sum_out_tmp[3][10];
        eta_sum[3][11]  = eta_sum_out_tmp[3][11];
        eta_sum[3][12]  = eta_sum_out_tmp[3][12];
        eta_sum[3][13]  = eta_sum_out_tmp[3][13];
        eta_sum[3][14]  = eta_sum_out_tmp[3][14];
        eta_sum[3][15]  = eta_sum_out_tmp[3][15];
        eta_sum[3][16]  = eta_sum_out_tmp[3][16];
        eta_sum[3][17]  = eta_sum_out_tmp[3][17];
        eta_sum[3][18]  = eta_sum_out_tmp[3][18];
        eta_sum[3][19]  = eta_sum_out_tmp[3][19];
        eta_sum[3][20]  = eta_sum_out_tmp[3][20];
        eta_sum[3][21]  = eta_sum_out_tmp[3][21];
        eta_sum[3][22]  = eta_sum_out_tmp[3][22];
        eta_sum[3][23]  = eta_sum_out_tmp[3][23];
        eta_sum[3][24]  = eta_sum_out_tmp[3][24];
        eta_sum[3][25]  = eta_sum_out_tmp[3][25];
        eta_sum[3][26]  = eta_sum_out_tmp[3][26];
        eta_sum[3][27]  = eta_sum_out_tmp[3][27];
        eta_sum[3][28]  = eta_sum_out_tmp[3][28];
        eta_sum[3][29]  = eta_sum_out_tmp[3][29];
        eta_sum[3][30]  = eta_sum_out_tmp[3][30];
        eta_sum[3][31]  = eta_sum_out_tmp[3][31];
        eta_sum[3][32]  = eta_sum_out_tmp[3][32];
        eta_sum[3][33]  = eta_sum_out_tmp[3][33];
        eta_sum[3][34]  = eta_sum_out_tmp[3][34];
        eta_sum[3][35]  = eta_sum_out_tmp[3][35];
        eta_sum[3][36]  = eta_sum_out_tmp[3][36];
        eta_sum[3][37]  = eta_sum_out_tmp[3][37];
        eta_sum[3][38]  = eta_sum_out_tmp[3][38];
        eta_sum[3][39]  = eta_sum_out_tmp[3][39];
        eta_sum[3][40]  = eta_sum_out_tmp[3][40];
        eta_sum[3][41]  = eta_sum_out_tmp[3][41];
    end
 
    1:begin 
        eta_sum[3][0]  = eta_sum_out_tmp[3][0];
        eta_sum[3][1]  = eta_sum_out_tmp[3][1];
        eta_sum[3][2]  = eta_sum_out_tmp[3][2];
        eta_sum[3][3]  = eta_sum_out_tmp[3][3];
        eta_sum[3][4]  = eta_sum_out_tmp[3][4];
        eta_sum[3][5]  = eta_sum_out_tmp[3][5];
        eta_sum[3][6]  = eta_sum_out_tmp[3][6];
        eta_sum[3][7]  = eta_sum_out_tmp[3][7];
        eta_sum[3][8]  = eta_sum_out_tmp[3][8];
        eta_sum[3][9]  = eta_sum_out_tmp[3][9];
        eta_sum[3][10]  = eta_sum_out_tmp[3][10];
        eta_sum[3][11]  = eta_sum_out_tmp[3][11];
        eta_sum[3][12]  = eta_sum_out_tmp[3][12];
        eta_sum[3][13]  = eta_sum_out_tmp[3][13];
        eta_sum[3][14]  = eta_sum_out_tmp[3][14];
        eta_sum[3][15]  = eta_sum_out_tmp[3][15];
        eta_sum[3][16]  = eta_sum_out_tmp[3][16];
        eta_sum[3][17]  = eta_sum_out_tmp[3][17];
        eta_sum[3][18]  = eta_sum_out_tmp[3][18];
        eta_sum[3][19]  = eta_sum_out_tmp[3][19];
        eta_sum[3][20]  = eta_sum_out_tmp[3][20];
        eta_sum[3][21]  = eta_sum_out_tmp[3][21];
        eta_sum[3][22]  = eta_sum_out_tmp[3][22];
        eta_sum[3][23]  = eta_sum_out_tmp[3][23];
        eta_sum[3][24]  = eta_sum_out_tmp[3][24];
        eta_sum[3][25]  = eta_sum_out_tmp[3][25];
        eta_sum[3][26]  = eta_sum_out_tmp[3][26];
        eta_sum[3][27]  = eta_sum_out_tmp[3][27];
        eta_sum[3][28]  = eta_sum_out_tmp[3][28];
        eta_sum[3][29]  = eta_sum_out_tmp[3][29];
        eta_sum[3][30]  = eta_sum_out_tmp[3][30];
        eta_sum[3][31]  = eta_sum_out_tmp[3][31];
        eta_sum[3][32]  = eta_sum_out_tmp[3][32];
        eta_sum[3][33]  = eta_sum_out_tmp[3][33];
        eta_sum[3][34]  = eta_sum_out_tmp[3][34];
        eta_sum[3][35]  = eta_sum_out_tmp[3][35];
        eta_sum[3][36]  = eta_sum_out_tmp[3][36];
        eta_sum[3][37]  = eta_sum_out_tmp[3][37];
        eta_sum[3][38]  = eta_sum_out_tmp[3][38];
        eta_sum[3][39]  = eta_sum_out_tmp[3][39];
        eta_sum[3][40]  = eta_sum_out_tmp[3][40];
        eta_sum[3][41]  = eta_sum_out_tmp[3][41];
    end
 
    2:begin 
        eta_sum[3][31]  = eta_sum_out_tmp[3][0];
        eta_sum[3][32]  = eta_sum_out_tmp[3][1];
        eta_sum[3][33]  = eta_sum_out_tmp[3][2];
        eta_sum[3][34]  = eta_sum_out_tmp[3][3];
        eta_sum[3][35]  = eta_sum_out_tmp[3][4];
        eta_sum[3][36]  = eta_sum_out_tmp[3][5];
        eta_sum[3][37]  = eta_sum_out_tmp[3][6];
        eta_sum[3][38]  = eta_sum_out_tmp[3][7];
        eta_sum[3][39]  = eta_sum_out_tmp[3][8];
        eta_sum[3][40]  = eta_sum_out_tmp[3][9];
        eta_sum[3][41]  = eta_sum_out_tmp[3][10];
        eta_sum[3][0]  = eta_sum_out_tmp[3][11];
        eta_sum[3][1]  = eta_sum_out_tmp[3][12];
        eta_sum[3][2]  = eta_sum_out_tmp[3][13];
        eta_sum[3][3]  = eta_sum_out_tmp[3][14];
        eta_sum[3][4]  = eta_sum_out_tmp[3][15];
        eta_sum[3][5]  = eta_sum_out_tmp[3][16];
        eta_sum[3][6]  = eta_sum_out_tmp[3][17];
        eta_sum[3][7]  = eta_sum_out_tmp[3][18];
        eta_sum[3][8]  = eta_sum_out_tmp[3][19];
        eta_sum[3][9]  = eta_sum_out_tmp[3][20];
        eta_sum[3][10]  = eta_sum_out_tmp[3][21];
        eta_sum[3][11]  = eta_sum_out_tmp[3][22];
        eta_sum[3][12]  = eta_sum_out_tmp[3][23];
        eta_sum[3][13]  = eta_sum_out_tmp[3][24];
        eta_sum[3][14]  = eta_sum_out_tmp[3][25];
        eta_sum[3][15]  = eta_sum_out_tmp[3][26];
        eta_sum[3][16]  = eta_sum_out_tmp[3][27];
        eta_sum[3][17]  = eta_sum_out_tmp[3][28];
        eta_sum[3][18]  = eta_sum_out_tmp[3][29];
        eta_sum[3][19]  = eta_sum_out_tmp[3][30];
        eta_sum[3][20]  = eta_sum_out_tmp[3][31];
        eta_sum[3][21]  = eta_sum_out_tmp[3][32];
        eta_sum[3][22]  = eta_sum_out_tmp[3][33];
        eta_sum[3][23]  = eta_sum_out_tmp[3][34];
        eta_sum[3][24]  = eta_sum_out_tmp[3][35];
        eta_sum[3][25]  = eta_sum_out_tmp[3][36];
        eta_sum[3][26]  = eta_sum_out_tmp[3][37];
        eta_sum[3][27]  = eta_sum_out_tmp[3][38];
        eta_sum[3][28]  = eta_sum_out_tmp[3][39];
        eta_sum[3][29]  = eta_sum_out_tmp[3][40];
        eta_sum[3][30]  = eta_sum_out_tmp[3][41];
    end
 
    3:begin 
        eta_sum[3][18]  = eta_sum_out_tmp[3][0];
        eta_sum[3][19]  = eta_sum_out_tmp[3][1];
        eta_sum[3][20]  = eta_sum_out_tmp[3][2];
        eta_sum[3][21]  = eta_sum_out_tmp[3][3];
        eta_sum[3][22]  = eta_sum_out_tmp[3][4];
        eta_sum[3][23]  = eta_sum_out_tmp[3][5];
        eta_sum[3][24]  = eta_sum_out_tmp[3][6];
        eta_sum[3][25]  = eta_sum_out_tmp[3][7];
        eta_sum[3][26]  = eta_sum_out_tmp[3][8];
        eta_sum[3][27]  = eta_sum_out_tmp[3][9];
        eta_sum[3][28]  = eta_sum_out_tmp[3][10];
        eta_sum[3][29]  = eta_sum_out_tmp[3][11];
        eta_sum[3][30]  = eta_sum_out_tmp[3][12];
        eta_sum[3][31]  = eta_sum_out_tmp[3][13];
        eta_sum[3][32]  = eta_sum_out_tmp[3][14];
        eta_sum[3][33]  = eta_sum_out_tmp[3][15];
        eta_sum[3][34]  = eta_sum_out_tmp[3][16];
        eta_sum[3][35]  = eta_sum_out_tmp[3][17];
        eta_sum[3][36]  = eta_sum_out_tmp[3][18];
        eta_sum[3][37]  = eta_sum_out_tmp[3][19];
        eta_sum[3][38]  = eta_sum_out_tmp[3][20];
        eta_sum[3][39]  = eta_sum_out_tmp[3][21];
        eta_sum[3][40]  = eta_sum_out_tmp[3][22];
        eta_sum[3][41]  = eta_sum_out_tmp[3][23];
        eta_sum[3][0]  = eta_sum_out_tmp[3][24];
        eta_sum[3][1]  = eta_sum_out_tmp[3][25];
        eta_sum[3][2]  = eta_sum_out_tmp[3][26];
        eta_sum[3][3]  = eta_sum_out_tmp[3][27];
        eta_sum[3][4]  = eta_sum_out_tmp[3][28];
        eta_sum[3][5]  = eta_sum_out_tmp[3][29];
        eta_sum[3][6]  = eta_sum_out_tmp[3][30];
        eta_sum[3][7]  = eta_sum_out_tmp[3][31];
        eta_sum[3][8]  = eta_sum_out_tmp[3][32];
        eta_sum[3][9]  = eta_sum_out_tmp[3][33];
        eta_sum[3][10]  = eta_sum_out_tmp[3][34];
        eta_sum[3][11]  = eta_sum_out_tmp[3][35];
        eta_sum[3][12]  = eta_sum_out_tmp[3][36];
        eta_sum[3][13]  = eta_sum_out_tmp[3][37];
        eta_sum[3][14]  = eta_sum_out_tmp[3][38];
        eta_sum[3][15]  = eta_sum_out_tmp[3][39];
        eta_sum[3][16]  = eta_sum_out_tmp[3][40];
        eta_sum[3][17]  = eta_sum_out_tmp[3][41];
    end
 
    4:begin 
        eta_sum[3][0]  = eta_sum_out_tmp[3][0];
        eta_sum[3][1]  = eta_sum_out_tmp[3][1];
        eta_sum[3][2]  = eta_sum_out_tmp[3][2];
        eta_sum[3][3]  = eta_sum_out_tmp[3][3];
        eta_sum[3][4]  = eta_sum_out_tmp[3][4];
        eta_sum[3][5]  = eta_sum_out_tmp[3][5];
        eta_sum[3][6]  = eta_sum_out_tmp[3][6];
        eta_sum[3][7]  = eta_sum_out_tmp[3][7];
        eta_sum[3][8]  = eta_sum_out_tmp[3][8];
        eta_sum[3][9]  = eta_sum_out_tmp[3][9];
        eta_sum[3][10]  = eta_sum_out_tmp[3][10];
        eta_sum[3][11]  = eta_sum_out_tmp[3][11];
        eta_sum[3][12]  = eta_sum_out_tmp[3][12];
        eta_sum[3][13]  = eta_sum_out_tmp[3][13];
        eta_sum[3][14]  = eta_sum_out_tmp[3][14];
        eta_sum[3][15]  = eta_sum_out_tmp[3][15];
        eta_sum[3][16]  = eta_sum_out_tmp[3][16];
        eta_sum[3][17]  = eta_sum_out_tmp[3][17];
        eta_sum[3][18]  = eta_sum_out_tmp[3][18];
        eta_sum[3][19]  = eta_sum_out_tmp[3][19];
        eta_sum[3][20]  = eta_sum_out_tmp[3][20];
        eta_sum[3][21]  = eta_sum_out_tmp[3][21];
        eta_sum[3][22]  = eta_sum_out_tmp[3][22];
        eta_sum[3][23]  = eta_sum_out_tmp[3][23];
        eta_sum[3][24]  = eta_sum_out_tmp[3][24];
        eta_sum[3][25]  = eta_sum_out_tmp[3][25];
        eta_sum[3][26]  = eta_sum_out_tmp[3][26];
        eta_sum[3][27]  = eta_sum_out_tmp[3][27];
        eta_sum[3][28]  = eta_sum_out_tmp[3][28];
        eta_sum[3][29]  = eta_sum_out_tmp[3][29];
        eta_sum[3][30]  = eta_sum_out_tmp[3][30];
        eta_sum[3][31]  = eta_sum_out_tmp[3][31];
        eta_sum[3][32]  = eta_sum_out_tmp[3][32];
        eta_sum[3][33]  = eta_sum_out_tmp[3][33];
        eta_sum[3][34]  = eta_sum_out_tmp[3][34];
        eta_sum[3][35]  = eta_sum_out_tmp[3][35];
        eta_sum[3][36]  = eta_sum_out_tmp[3][36];
        eta_sum[3][37]  = eta_sum_out_tmp[3][37];
        eta_sum[3][38]  = eta_sum_out_tmp[3][38];
        eta_sum[3][39]  = eta_sum_out_tmp[3][39];
        eta_sum[3][40]  = eta_sum_out_tmp[3][40];
        eta_sum[3][41]  = eta_sum_out_tmp[3][41];
    end
 
    5:begin 
        eta_sum[3][0]  = eta_sum_out_tmp[3][0];
        eta_sum[3][1]  = eta_sum_out_tmp[3][1];
        eta_sum[3][2]  = eta_sum_out_tmp[3][2];
        eta_sum[3][3]  = eta_sum_out_tmp[3][3];
        eta_sum[3][4]  = eta_sum_out_tmp[3][4];
        eta_sum[3][5]  = eta_sum_out_tmp[3][5];
        eta_sum[3][6]  = eta_sum_out_tmp[3][6];
        eta_sum[3][7]  = eta_sum_out_tmp[3][7];
        eta_sum[3][8]  = eta_sum_out_tmp[3][8];
        eta_sum[3][9]  = eta_sum_out_tmp[3][9];
        eta_sum[3][10]  = eta_sum_out_tmp[3][10];
        eta_sum[3][11]  = eta_sum_out_tmp[3][11];
        eta_sum[3][12]  = eta_sum_out_tmp[3][12];
        eta_sum[3][13]  = eta_sum_out_tmp[3][13];
        eta_sum[3][14]  = eta_sum_out_tmp[3][14];
        eta_sum[3][15]  = eta_sum_out_tmp[3][15];
        eta_sum[3][16]  = eta_sum_out_tmp[3][16];
        eta_sum[3][17]  = eta_sum_out_tmp[3][17];
        eta_sum[3][18]  = eta_sum_out_tmp[3][18];
        eta_sum[3][19]  = eta_sum_out_tmp[3][19];
        eta_sum[3][20]  = eta_sum_out_tmp[3][20];
        eta_sum[3][21]  = eta_sum_out_tmp[3][21];
        eta_sum[3][22]  = eta_sum_out_tmp[3][22];
        eta_sum[3][23]  = eta_sum_out_tmp[3][23];
        eta_sum[3][24]  = eta_sum_out_tmp[3][24];
        eta_sum[3][25]  = eta_sum_out_tmp[3][25];
        eta_sum[3][26]  = eta_sum_out_tmp[3][26];
        eta_sum[3][27]  = eta_sum_out_tmp[3][27];
        eta_sum[3][28]  = eta_sum_out_tmp[3][28];
        eta_sum[3][29]  = eta_sum_out_tmp[3][29];
        eta_sum[3][30]  = eta_sum_out_tmp[3][30];
        eta_sum[3][31]  = eta_sum_out_tmp[3][31];
        eta_sum[3][32]  = eta_sum_out_tmp[3][32];
        eta_sum[3][33]  = eta_sum_out_tmp[3][33];
        eta_sum[3][34]  = eta_sum_out_tmp[3][34];
        eta_sum[3][35]  = eta_sum_out_tmp[3][35];
        eta_sum[3][36]  = eta_sum_out_tmp[3][36];
        eta_sum[3][37]  = eta_sum_out_tmp[3][37];
        eta_sum[3][38]  = eta_sum_out_tmp[3][38];
        eta_sum[3][39]  = eta_sum_out_tmp[3][39];
        eta_sum[3][40]  = eta_sum_out_tmp[3][40];
        eta_sum[3][41]  = eta_sum_out_tmp[3][41];
    end
 
    6:begin 
        eta_sum[3][23]  = eta_sum_out_tmp[3][0];
        eta_sum[3][24]  = eta_sum_out_tmp[3][1];
        eta_sum[3][25]  = eta_sum_out_tmp[3][2];
        eta_sum[3][26]  = eta_sum_out_tmp[3][3];
        eta_sum[3][27]  = eta_sum_out_tmp[3][4];
        eta_sum[3][28]  = eta_sum_out_tmp[3][5];
        eta_sum[3][29]  = eta_sum_out_tmp[3][6];
        eta_sum[3][30]  = eta_sum_out_tmp[3][7];
        eta_sum[3][31]  = eta_sum_out_tmp[3][8];
        eta_sum[3][32]  = eta_sum_out_tmp[3][9];
        eta_sum[3][33]  = eta_sum_out_tmp[3][10];
        eta_sum[3][34]  = eta_sum_out_tmp[3][11];
        eta_sum[3][35]  = eta_sum_out_tmp[3][12];
        eta_sum[3][36]  = eta_sum_out_tmp[3][13];
        eta_sum[3][37]  = eta_sum_out_tmp[3][14];
        eta_sum[3][38]  = eta_sum_out_tmp[3][15];
        eta_sum[3][39]  = eta_sum_out_tmp[3][16];
        eta_sum[3][40]  = eta_sum_out_tmp[3][17];
        eta_sum[3][41]  = eta_sum_out_tmp[3][18];
        eta_sum[3][0]  = eta_sum_out_tmp[3][19];
        eta_sum[3][1]  = eta_sum_out_tmp[3][20];
        eta_sum[3][2]  = eta_sum_out_tmp[3][21];
        eta_sum[3][3]  = eta_sum_out_tmp[3][22];
        eta_sum[3][4]  = eta_sum_out_tmp[3][23];
        eta_sum[3][5]  = eta_sum_out_tmp[3][24];
        eta_sum[3][6]  = eta_sum_out_tmp[3][25];
        eta_sum[3][7]  = eta_sum_out_tmp[3][26];
        eta_sum[3][8]  = eta_sum_out_tmp[3][27];
        eta_sum[3][9]  = eta_sum_out_tmp[3][28];
        eta_sum[3][10]  = eta_sum_out_tmp[3][29];
        eta_sum[3][11]  = eta_sum_out_tmp[3][30];
        eta_sum[3][12]  = eta_sum_out_tmp[3][31];
        eta_sum[3][13]  = eta_sum_out_tmp[3][32];
        eta_sum[3][14]  = eta_sum_out_tmp[3][33];
        eta_sum[3][15]  = eta_sum_out_tmp[3][34];
        eta_sum[3][16]  = eta_sum_out_tmp[3][35];
        eta_sum[3][17]  = eta_sum_out_tmp[3][36];
        eta_sum[3][18]  = eta_sum_out_tmp[3][37];
        eta_sum[3][19]  = eta_sum_out_tmp[3][38];
        eta_sum[3][20]  = eta_sum_out_tmp[3][39];
        eta_sum[3][21]  = eta_sum_out_tmp[3][40];
        eta_sum[3][22]  = eta_sum_out_tmp[3][41];
    end
 
    7:begin 
        eta_sum[3][34]  = eta_sum_out_tmp[3][0];
        eta_sum[3][35]  = eta_sum_out_tmp[3][1];
        eta_sum[3][36]  = eta_sum_out_tmp[3][2];
        eta_sum[3][37]  = eta_sum_out_tmp[3][3];
        eta_sum[3][38]  = eta_sum_out_tmp[3][4];
        eta_sum[3][39]  = eta_sum_out_tmp[3][5];
        eta_sum[3][40]  = eta_sum_out_tmp[3][6];
        eta_sum[3][41]  = eta_sum_out_tmp[3][7];
        eta_sum[3][0]  = eta_sum_out_tmp[3][8];
        eta_sum[3][1]  = eta_sum_out_tmp[3][9];
        eta_sum[3][2]  = eta_sum_out_tmp[3][10];
        eta_sum[3][3]  = eta_sum_out_tmp[3][11];
        eta_sum[3][4]  = eta_sum_out_tmp[3][12];
        eta_sum[3][5]  = eta_sum_out_tmp[3][13];
        eta_sum[3][6]  = eta_sum_out_tmp[3][14];
        eta_sum[3][7]  = eta_sum_out_tmp[3][15];
        eta_sum[3][8]  = eta_sum_out_tmp[3][16];
        eta_sum[3][9]  = eta_sum_out_tmp[3][17];
        eta_sum[3][10]  = eta_sum_out_tmp[3][18];
        eta_sum[3][11]  = eta_sum_out_tmp[3][19];
        eta_sum[3][12]  = eta_sum_out_tmp[3][20];
        eta_sum[3][13]  = eta_sum_out_tmp[3][21];
        eta_sum[3][14]  = eta_sum_out_tmp[3][22];
        eta_sum[3][15]  = eta_sum_out_tmp[3][23];
        eta_sum[3][16]  = eta_sum_out_tmp[3][24];
        eta_sum[3][17]  = eta_sum_out_tmp[3][25];
        eta_sum[3][18]  = eta_sum_out_tmp[3][26];
        eta_sum[3][19]  = eta_sum_out_tmp[3][27];
        eta_sum[3][20]  = eta_sum_out_tmp[3][28];
        eta_sum[3][21]  = eta_sum_out_tmp[3][29];
        eta_sum[3][22]  = eta_sum_out_tmp[3][30];
        eta_sum[3][23]  = eta_sum_out_tmp[3][31];
        eta_sum[3][24]  = eta_sum_out_tmp[3][32];
        eta_sum[3][25]  = eta_sum_out_tmp[3][33];
        eta_sum[3][26]  = eta_sum_out_tmp[3][34];
        eta_sum[3][27]  = eta_sum_out_tmp[3][35];
        eta_sum[3][28]  = eta_sum_out_tmp[3][36];
        eta_sum[3][29]  = eta_sum_out_tmp[3][37];
        eta_sum[3][30]  = eta_sum_out_tmp[3][38];
        eta_sum[3][31]  = eta_sum_out_tmp[3][39];
        eta_sum[3][32]  = eta_sum_out_tmp[3][40];
        eta_sum[3][33]  = eta_sum_out_tmp[3][41];
    end
 
endcase
end

if (chk_n_output_valid[0] & active_cols[4]) begin
case (curr_layer)
    0:begin 
        eta_sum[4][13]  = eta_sum_out_tmp[4][0];
        eta_sum[4][14]  = eta_sum_out_tmp[4][1];
        eta_sum[4][15]  = eta_sum_out_tmp[4][2];
        eta_sum[4][16]  = eta_sum_out_tmp[4][3];
        eta_sum[4][17]  = eta_sum_out_tmp[4][4];
        eta_sum[4][18]  = eta_sum_out_tmp[4][5];
        eta_sum[4][19]  = eta_sum_out_tmp[4][6];
        eta_sum[4][20]  = eta_sum_out_tmp[4][7];
        eta_sum[4][21]  = eta_sum_out_tmp[4][8];
        eta_sum[4][22]  = eta_sum_out_tmp[4][9];
        eta_sum[4][23]  = eta_sum_out_tmp[4][10];
        eta_sum[4][24]  = eta_sum_out_tmp[4][11];
        eta_sum[4][25]  = eta_sum_out_tmp[4][12];
        eta_sum[4][26]  = eta_sum_out_tmp[4][13];
        eta_sum[4][27]  = eta_sum_out_tmp[4][14];
        eta_sum[4][28]  = eta_sum_out_tmp[4][15];
        eta_sum[4][29]  = eta_sum_out_tmp[4][16];
        eta_sum[4][30]  = eta_sum_out_tmp[4][17];
        eta_sum[4][31]  = eta_sum_out_tmp[4][18];
        eta_sum[4][32]  = eta_sum_out_tmp[4][19];
        eta_sum[4][33]  = eta_sum_out_tmp[4][20];
        eta_sum[4][34]  = eta_sum_out_tmp[4][21];
        eta_sum[4][35]  = eta_sum_out_tmp[4][22];
        eta_sum[4][36]  = eta_sum_out_tmp[4][23];
        eta_sum[4][37]  = eta_sum_out_tmp[4][24];
        eta_sum[4][38]  = eta_sum_out_tmp[4][25];
        eta_sum[4][39]  = eta_sum_out_tmp[4][26];
        eta_sum[4][40]  = eta_sum_out_tmp[4][27];
        eta_sum[4][41]  = eta_sum_out_tmp[4][28];
        eta_sum[4][0]  = eta_sum_out_tmp[4][29];
        eta_sum[4][1]  = eta_sum_out_tmp[4][30];
        eta_sum[4][2]  = eta_sum_out_tmp[4][31];
        eta_sum[4][3]  = eta_sum_out_tmp[4][32];
        eta_sum[4][4]  = eta_sum_out_tmp[4][33];
        eta_sum[4][5]  = eta_sum_out_tmp[4][34];
        eta_sum[4][6]  = eta_sum_out_tmp[4][35];
        eta_sum[4][7]  = eta_sum_out_tmp[4][36];
        eta_sum[4][8]  = eta_sum_out_tmp[4][37];
        eta_sum[4][9]  = eta_sum_out_tmp[4][38];
        eta_sum[4][10]  = eta_sum_out_tmp[4][39];
        eta_sum[4][11]  = eta_sum_out_tmp[4][40];
        eta_sum[4][12]  = eta_sum_out_tmp[4][41];
    end
 
    1:begin 
        eta_sum[4][27]  = eta_sum_out_tmp[4][0];
        eta_sum[4][28]  = eta_sum_out_tmp[4][1];
        eta_sum[4][29]  = eta_sum_out_tmp[4][2];
        eta_sum[4][30]  = eta_sum_out_tmp[4][3];
        eta_sum[4][31]  = eta_sum_out_tmp[4][4];
        eta_sum[4][32]  = eta_sum_out_tmp[4][5];
        eta_sum[4][33]  = eta_sum_out_tmp[4][6];
        eta_sum[4][34]  = eta_sum_out_tmp[4][7];
        eta_sum[4][35]  = eta_sum_out_tmp[4][8];
        eta_sum[4][36]  = eta_sum_out_tmp[4][9];
        eta_sum[4][37]  = eta_sum_out_tmp[4][10];
        eta_sum[4][38]  = eta_sum_out_tmp[4][11];
        eta_sum[4][39]  = eta_sum_out_tmp[4][12];
        eta_sum[4][40]  = eta_sum_out_tmp[4][13];
        eta_sum[4][41]  = eta_sum_out_tmp[4][14];
        eta_sum[4][0]  = eta_sum_out_tmp[4][15];
        eta_sum[4][1]  = eta_sum_out_tmp[4][16];
        eta_sum[4][2]  = eta_sum_out_tmp[4][17];
        eta_sum[4][3]  = eta_sum_out_tmp[4][18];
        eta_sum[4][4]  = eta_sum_out_tmp[4][19];
        eta_sum[4][5]  = eta_sum_out_tmp[4][20];
        eta_sum[4][6]  = eta_sum_out_tmp[4][21];
        eta_sum[4][7]  = eta_sum_out_tmp[4][22];
        eta_sum[4][8]  = eta_sum_out_tmp[4][23];
        eta_sum[4][9]  = eta_sum_out_tmp[4][24];
        eta_sum[4][10]  = eta_sum_out_tmp[4][25];
        eta_sum[4][11]  = eta_sum_out_tmp[4][26];
        eta_sum[4][12]  = eta_sum_out_tmp[4][27];
        eta_sum[4][13]  = eta_sum_out_tmp[4][28];
        eta_sum[4][14]  = eta_sum_out_tmp[4][29];
        eta_sum[4][15]  = eta_sum_out_tmp[4][30];
        eta_sum[4][16]  = eta_sum_out_tmp[4][31];
        eta_sum[4][17]  = eta_sum_out_tmp[4][32];
        eta_sum[4][18]  = eta_sum_out_tmp[4][33];
        eta_sum[4][19]  = eta_sum_out_tmp[4][34];
        eta_sum[4][20]  = eta_sum_out_tmp[4][35];
        eta_sum[4][21]  = eta_sum_out_tmp[4][36];
        eta_sum[4][22]  = eta_sum_out_tmp[4][37];
        eta_sum[4][23]  = eta_sum_out_tmp[4][38];
        eta_sum[4][24]  = eta_sum_out_tmp[4][39];
        eta_sum[4][25]  = eta_sum_out_tmp[4][40];
        eta_sum[4][26]  = eta_sum_out_tmp[4][41];
    end
 
    2:begin 
        eta_sum[4][0]  = eta_sum_out_tmp[4][0];
        eta_sum[4][1]  = eta_sum_out_tmp[4][1];
        eta_sum[4][2]  = eta_sum_out_tmp[4][2];
        eta_sum[4][3]  = eta_sum_out_tmp[4][3];
        eta_sum[4][4]  = eta_sum_out_tmp[4][4];
        eta_sum[4][5]  = eta_sum_out_tmp[4][5];
        eta_sum[4][6]  = eta_sum_out_tmp[4][6];
        eta_sum[4][7]  = eta_sum_out_tmp[4][7];
        eta_sum[4][8]  = eta_sum_out_tmp[4][8];
        eta_sum[4][9]  = eta_sum_out_tmp[4][9];
        eta_sum[4][10]  = eta_sum_out_tmp[4][10];
        eta_sum[4][11]  = eta_sum_out_tmp[4][11];
        eta_sum[4][12]  = eta_sum_out_tmp[4][12];
        eta_sum[4][13]  = eta_sum_out_tmp[4][13];
        eta_sum[4][14]  = eta_sum_out_tmp[4][14];
        eta_sum[4][15]  = eta_sum_out_tmp[4][15];
        eta_sum[4][16]  = eta_sum_out_tmp[4][16];
        eta_sum[4][17]  = eta_sum_out_tmp[4][17];
        eta_sum[4][18]  = eta_sum_out_tmp[4][18];
        eta_sum[4][19]  = eta_sum_out_tmp[4][19];
        eta_sum[4][20]  = eta_sum_out_tmp[4][20];
        eta_sum[4][21]  = eta_sum_out_tmp[4][21];
        eta_sum[4][22]  = eta_sum_out_tmp[4][22];
        eta_sum[4][23]  = eta_sum_out_tmp[4][23];
        eta_sum[4][24]  = eta_sum_out_tmp[4][24];
        eta_sum[4][25]  = eta_sum_out_tmp[4][25];
        eta_sum[4][26]  = eta_sum_out_tmp[4][26];
        eta_sum[4][27]  = eta_sum_out_tmp[4][27];
        eta_sum[4][28]  = eta_sum_out_tmp[4][28];
        eta_sum[4][29]  = eta_sum_out_tmp[4][29];
        eta_sum[4][30]  = eta_sum_out_tmp[4][30];
        eta_sum[4][31]  = eta_sum_out_tmp[4][31];
        eta_sum[4][32]  = eta_sum_out_tmp[4][32];
        eta_sum[4][33]  = eta_sum_out_tmp[4][33];
        eta_sum[4][34]  = eta_sum_out_tmp[4][34];
        eta_sum[4][35]  = eta_sum_out_tmp[4][35];
        eta_sum[4][36]  = eta_sum_out_tmp[4][36];
        eta_sum[4][37]  = eta_sum_out_tmp[4][37];
        eta_sum[4][38]  = eta_sum_out_tmp[4][38];
        eta_sum[4][39]  = eta_sum_out_tmp[4][39];
        eta_sum[4][40]  = eta_sum_out_tmp[4][40];
        eta_sum[4][41]  = eta_sum_out_tmp[4][41];
    end
 
    3:begin 
        eta_sum[4][0]  = eta_sum_out_tmp[4][0];
        eta_sum[4][1]  = eta_sum_out_tmp[4][1];
        eta_sum[4][2]  = eta_sum_out_tmp[4][2];
        eta_sum[4][3]  = eta_sum_out_tmp[4][3];
        eta_sum[4][4]  = eta_sum_out_tmp[4][4];
        eta_sum[4][5]  = eta_sum_out_tmp[4][5];
        eta_sum[4][6]  = eta_sum_out_tmp[4][6];
        eta_sum[4][7]  = eta_sum_out_tmp[4][7];
        eta_sum[4][8]  = eta_sum_out_tmp[4][8];
        eta_sum[4][9]  = eta_sum_out_tmp[4][9];
        eta_sum[4][10]  = eta_sum_out_tmp[4][10];
        eta_sum[4][11]  = eta_sum_out_tmp[4][11];
        eta_sum[4][12]  = eta_sum_out_tmp[4][12];
        eta_sum[4][13]  = eta_sum_out_tmp[4][13];
        eta_sum[4][14]  = eta_sum_out_tmp[4][14];
        eta_sum[4][15]  = eta_sum_out_tmp[4][15];
        eta_sum[4][16]  = eta_sum_out_tmp[4][16];
        eta_sum[4][17]  = eta_sum_out_tmp[4][17];
        eta_sum[4][18]  = eta_sum_out_tmp[4][18];
        eta_sum[4][19]  = eta_sum_out_tmp[4][19];
        eta_sum[4][20]  = eta_sum_out_tmp[4][20];
        eta_sum[4][21]  = eta_sum_out_tmp[4][21];
        eta_sum[4][22]  = eta_sum_out_tmp[4][22];
        eta_sum[4][23]  = eta_sum_out_tmp[4][23];
        eta_sum[4][24]  = eta_sum_out_tmp[4][24];
        eta_sum[4][25]  = eta_sum_out_tmp[4][25];
        eta_sum[4][26]  = eta_sum_out_tmp[4][26];
        eta_sum[4][27]  = eta_sum_out_tmp[4][27];
        eta_sum[4][28]  = eta_sum_out_tmp[4][28];
        eta_sum[4][29]  = eta_sum_out_tmp[4][29];
        eta_sum[4][30]  = eta_sum_out_tmp[4][30];
        eta_sum[4][31]  = eta_sum_out_tmp[4][31];
        eta_sum[4][32]  = eta_sum_out_tmp[4][32];
        eta_sum[4][33]  = eta_sum_out_tmp[4][33];
        eta_sum[4][34]  = eta_sum_out_tmp[4][34];
        eta_sum[4][35]  = eta_sum_out_tmp[4][35];
        eta_sum[4][36]  = eta_sum_out_tmp[4][36];
        eta_sum[4][37]  = eta_sum_out_tmp[4][37];
        eta_sum[4][38]  = eta_sum_out_tmp[4][38];
        eta_sum[4][39]  = eta_sum_out_tmp[4][39];
        eta_sum[4][40]  = eta_sum_out_tmp[4][40];
        eta_sum[4][41]  = eta_sum_out_tmp[4][41];
    end
 
    4:begin 
        eta_sum[4][40]  = eta_sum_out_tmp[4][0];
        eta_sum[4][41]  = eta_sum_out_tmp[4][1];
        eta_sum[4][0]  = eta_sum_out_tmp[4][2];
        eta_sum[4][1]  = eta_sum_out_tmp[4][3];
        eta_sum[4][2]  = eta_sum_out_tmp[4][4];
        eta_sum[4][3]  = eta_sum_out_tmp[4][5];
        eta_sum[4][4]  = eta_sum_out_tmp[4][6];
        eta_sum[4][5]  = eta_sum_out_tmp[4][7];
        eta_sum[4][6]  = eta_sum_out_tmp[4][8];
        eta_sum[4][7]  = eta_sum_out_tmp[4][9];
        eta_sum[4][8]  = eta_sum_out_tmp[4][10];
        eta_sum[4][9]  = eta_sum_out_tmp[4][11];
        eta_sum[4][10]  = eta_sum_out_tmp[4][12];
        eta_sum[4][11]  = eta_sum_out_tmp[4][13];
        eta_sum[4][12]  = eta_sum_out_tmp[4][14];
        eta_sum[4][13]  = eta_sum_out_tmp[4][15];
        eta_sum[4][14]  = eta_sum_out_tmp[4][16];
        eta_sum[4][15]  = eta_sum_out_tmp[4][17];
        eta_sum[4][16]  = eta_sum_out_tmp[4][18];
        eta_sum[4][17]  = eta_sum_out_tmp[4][19];
        eta_sum[4][18]  = eta_sum_out_tmp[4][20];
        eta_sum[4][19]  = eta_sum_out_tmp[4][21];
        eta_sum[4][20]  = eta_sum_out_tmp[4][22];
        eta_sum[4][21]  = eta_sum_out_tmp[4][23];
        eta_sum[4][22]  = eta_sum_out_tmp[4][24];
        eta_sum[4][23]  = eta_sum_out_tmp[4][25];
        eta_sum[4][24]  = eta_sum_out_tmp[4][26];
        eta_sum[4][25]  = eta_sum_out_tmp[4][27];
        eta_sum[4][26]  = eta_sum_out_tmp[4][28];
        eta_sum[4][27]  = eta_sum_out_tmp[4][29];
        eta_sum[4][28]  = eta_sum_out_tmp[4][30];
        eta_sum[4][29]  = eta_sum_out_tmp[4][31];
        eta_sum[4][30]  = eta_sum_out_tmp[4][32];
        eta_sum[4][31]  = eta_sum_out_tmp[4][33];
        eta_sum[4][32]  = eta_sum_out_tmp[4][34];
        eta_sum[4][33]  = eta_sum_out_tmp[4][35];
        eta_sum[4][34]  = eta_sum_out_tmp[4][36];
        eta_sum[4][35]  = eta_sum_out_tmp[4][37];
        eta_sum[4][36]  = eta_sum_out_tmp[4][38];
        eta_sum[4][37]  = eta_sum_out_tmp[4][39];
        eta_sum[4][38]  = eta_sum_out_tmp[4][40];
        eta_sum[4][39]  = eta_sum_out_tmp[4][41];
    end
 
    5:begin 
        eta_sum[4][0]  = eta_sum_out_tmp[4][0];
        eta_sum[4][1]  = eta_sum_out_tmp[4][1];
        eta_sum[4][2]  = eta_sum_out_tmp[4][2];
        eta_sum[4][3]  = eta_sum_out_tmp[4][3];
        eta_sum[4][4]  = eta_sum_out_tmp[4][4];
        eta_sum[4][5]  = eta_sum_out_tmp[4][5];
        eta_sum[4][6]  = eta_sum_out_tmp[4][6];
        eta_sum[4][7]  = eta_sum_out_tmp[4][7];
        eta_sum[4][8]  = eta_sum_out_tmp[4][8];
        eta_sum[4][9]  = eta_sum_out_tmp[4][9];
        eta_sum[4][10]  = eta_sum_out_tmp[4][10];
        eta_sum[4][11]  = eta_sum_out_tmp[4][11];
        eta_sum[4][12]  = eta_sum_out_tmp[4][12];
        eta_sum[4][13]  = eta_sum_out_tmp[4][13];
        eta_sum[4][14]  = eta_sum_out_tmp[4][14];
        eta_sum[4][15]  = eta_sum_out_tmp[4][15];
        eta_sum[4][16]  = eta_sum_out_tmp[4][16];
        eta_sum[4][17]  = eta_sum_out_tmp[4][17];
        eta_sum[4][18]  = eta_sum_out_tmp[4][18];
        eta_sum[4][19]  = eta_sum_out_tmp[4][19];
        eta_sum[4][20]  = eta_sum_out_tmp[4][20];
        eta_sum[4][21]  = eta_sum_out_tmp[4][21];
        eta_sum[4][22]  = eta_sum_out_tmp[4][22];
        eta_sum[4][23]  = eta_sum_out_tmp[4][23];
        eta_sum[4][24]  = eta_sum_out_tmp[4][24];
        eta_sum[4][25]  = eta_sum_out_tmp[4][25];
        eta_sum[4][26]  = eta_sum_out_tmp[4][26];
        eta_sum[4][27]  = eta_sum_out_tmp[4][27];
        eta_sum[4][28]  = eta_sum_out_tmp[4][28];
        eta_sum[4][29]  = eta_sum_out_tmp[4][29];
        eta_sum[4][30]  = eta_sum_out_tmp[4][30];
        eta_sum[4][31]  = eta_sum_out_tmp[4][31];
        eta_sum[4][32]  = eta_sum_out_tmp[4][32];
        eta_sum[4][33]  = eta_sum_out_tmp[4][33];
        eta_sum[4][34]  = eta_sum_out_tmp[4][34];
        eta_sum[4][35]  = eta_sum_out_tmp[4][35];
        eta_sum[4][36]  = eta_sum_out_tmp[4][36];
        eta_sum[4][37]  = eta_sum_out_tmp[4][37];
        eta_sum[4][38]  = eta_sum_out_tmp[4][38];
        eta_sum[4][39]  = eta_sum_out_tmp[4][39];
        eta_sum[4][40]  = eta_sum_out_tmp[4][40];
        eta_sum[4][41]  = eta_sum_out_tmp[4][41];
    end
 
    6:begin 
        eta_sum[4][0]  = eta_sum_out_tmp[4][0];
        eta_sum[4][1]  = eta_sum_out_tmp[4][1];
        eta_sum[4][2]  = eta_sum_out_tmp[4][2];
        eta_sum[4][3]  = eta_sum_out_tmp[4][3];
        eta_sum[4][4]  = eta_sum_out_tmp[4][4];
        eta_sum[4][5]  = eta_sum_out_tmp[4][5];
        eta_sum[4][6]  = eta_sum_out_tmp[4][6];
        eta_sum[4][7]  = eta_sum_out_tmp[4][7];
        eta_sum[4][8]  = eta_sum_out_tmp[4][8];
        eta_sum[4][9]  = eta_sum_out_tmp[4][9];
        eta_sum[4][10]  = eta_sum_out_tmp[4][10];
        eta_sum[4][11]  = eta_sum_out_tmp[4][11];
        eta_sum[4][12]  = eta_sum_out_tmp[4][12];
        eta_sum[4][13]  = eta_sum_out_tmp[4][13];
        eta_sum[4][14]  = eta_sum_out_tmp[4][14];
        eta_sum[4][15]  = eta_sum_out_tmp[4][15];
        eta_sum[4][16]  = eta_sum_out_tmp[4][16];
        eta_sum[4][17]  = eta_sum_out_tmp[4][17];
        eta_sum[4][18]  = eta_sum_out_tmp[4][18];
        eta_sum[4][19]  = eta_sum_out_tmp[4][19];
        eta_sum[4][20]  = eta_sum_out_tmp[4][20];
        eta_sum[4][21]  = eta_sum_out_tmp[4][21];
        eta_sum[4][22]  = eta_sum_out_tmp[4][22];
        eta_sum[4][23]  = eta_sum_out_tmp[4][23];
        eta_sum[4][24]  = eta_sum_out_tmp[4][24];
        eta_sum[4][25]  = eta_sum_out_tmp[4][25];
        eta_sum[4][26]  = eta_sum_out_tmp[4][26];
        eta_sum[4][27]  = eta_sum_out_tmp[4][27];
        eta_sum[4][28]  = eta_sum_out_tmp[4][28];
        eta_sum[4][29]  = eta_sum_out_tmp[4][29];
        eta_sum[4][30]  = eta_sum_out_tmp[4][30];
        eta_sum[4][31]  = eta_sum_out_tmp[4][31];
        eta_sum[4][32]  = eta_sum_out_tmp[4][32];
        eta_sum[4][33]  = eta_sum_out_tmp[4][33];
        eta_sum[4][34]  = eta_sum_out_tmp[4][34];
        eta_sum[4][35]  = eta_sum_out_tmp[4][35];
        eta_sum[4][36]  = eta_sum_out_tmp[4][36];
        eta_sum[4][37]  = eta_sum_out_tmp[4][37];
        eta_sum[4][38]  = eta_sum_out_tmp[4][38];
        eta_sum[4][39]  = eta_sum_out_tmp[4][39];
        eta_sum[4][40]  = eta_sum_out_tmp[4][40];
        eta_sum[4][41]  = eta_sum_out_tmp[4][41];
    end
 
    7:begin 
        eta_sum[4][31]  = eta_sum_out_tmp[4][0];
        eta_sum[4][32]  = eta_sum_out_tmp[4][1];
        eta_sum[4][33]  = eta_sum_out_tmp[4][2];
        eta_sum[4][34]  = eta_sum_out_tmp[4][3];
        eta_sum[4][35]  = eta_sum_out_tmp[4][4];
        eta_sum[4][36]  = eta_sum_out_tmp[4][5];
        eta_sum[4][37]  = eta_sum_out_tmp[4][6];
        eta_sum[4][38]  = eta_sum_out_tmp[4][7];
        eta_sum[4][39]  = eta_sum_out_tmp[4][8];
        eta_sum[4][40]  = eta_sum_out_tmp[4][9];
        eta_sum[4][41]  = eta_sum_out_tmp[4][10];
        eta_sum[4][0]  = eta_sum_out_tmp[4][11];
        eta_sum[4][1]  = eta_sum_out_tmp[4][12];
        eta_sum[4][2]  = eta_sum_out_tmp[4][13];
        eta_sum[4][3]  = eta_sum_out_tmp[4][14];
        eta_sum[4][4]  = eta_sum_out_tmp[4][15];
        eta_sum[4][5]  = eta_sum_out_tmp[4][16];
        eta_sum[4][6]  = eta_sum_out_tmp[4][17];
        eta_sum[4][7]  = eta_sum_out_tmp[4][18];
        eta_sum[4][8]  = eta_sum_out_tmp[4][19];
        eta_sum[4][9]  = eta_sum_out_tmp[4][20];
        eta_sum[4][10]  = eta_sum_out_tmp[4][21];
        eta_sum[4][11]  = eta_sum_out_tmp[4][22];
        eta_sum[4][12]  = eta_sum_out_tmp[4][23];
        eta_sum[4][13]  = eta_sum_out_tmp[4][24];
        eta_sum[4][14]  = eta_sum_out_tmp[4][25];
        eta_sum[4][15]  = eta_sum_out_tmp[4][26];
        eta_sum[4][16]  = eta_sum_out_tmp[4][27];
        eta_sum[4][17]  = eta_sum_out_tmp[4][28];
        eta_sum[4][18]  = eta_sum_out_tmp[4][29];
        eta_sum[4][19]  = eta_sum_out_tmp[4][30];
        eta_sum[4][20]  = eta_sum_out_tmp[4][31];
        eta_sum[4][21]  = eta_sum_out_tmp[4][32];
        eta_sum[4][22]  = eta_sum_out_tmp[4][33];
        eta_sum[4][23]  = eta_sum_out_tmp[4][34];
        eta_sum[4][24]  = eta_sum_out_tmp[4][35];
        eta_sum[4][25]  = eta_sum_out_tmp[4][36];
        eta_sum[4][26]  = eta_sum_out_tmp[4][37];
        eta_sum[4][27]  = eta_sum_out_tmp[4][38];
        eta_sum[4][28]  = eta_sum_out_tmp[4][39];
        eta_sum[4][29]  = eta_sum_out_tmp[4][40];
        eta_sum[4][30]  = eta_sum_out_tmp[4][41];
    end
 
endcase
end

if (chk_n_output_valid[0] & active_cols[5]) begin
case (curr_layer)
    0:begin 
        eta_sum[5][0]  = eta_sum_out_tmp[5][0];
        eta_sum[5][1]  = eta_sum_out_tmp[5][1];
        eta_sum[5][2]  = eta_sum_out_tmp[5][2];
        eta_sum[5][3]  = eta_sum_out_tmp[5][3];
        eta_sum[5][4]  = eta_sum_out_tmp[5][4];
        eta_sum[5][5]  = eta_sum_out_tmp[5][5];
        eta_sum[5][6]  = eta_sum_out_tmp[5][6];
        eta_sum[5][7]  = eta_sum_out_tmp[5][7];
        eta_sum[5][8]  = eta_sum_out_tmp[5][8];
        eta_sum[5][9]  = eta_sum_out_tmp[5][9];
        eta_sum[5][10]  = eta_sum_out_tmp[5][10];
        eta_sum[5][11]  = eta_sum_out_tmp[5][11];
        eta_sum[5][12]  = eta_sum_out_tmp[5][12];
        eta_sum[5][13]  = eta_sum_out_tmp[5][13];
        eta_sum[5][14]  = eta_sum_out_tmp[5][14];
        eta_sum[5][15]  = eta_sum_out_tmp[5][15];
        eta_sum[5][16]  = eta_sum_out_tmp[5][16];
        eta_sum[5][17]  = eta_sum_out_tmp[5][17];
        eta_sum[5][18]  = eta_sum_out_tmp[5][18];
        eta_sum[5][19]  = eta_sum_out_tmp[5][19];
        eta_sum[5][20]  = eta_sum_out_tmp[5][20];
        eta_sum[5][21]  = eta_sum_out_tmp[5][21];
        eta_sum[5][22]  = eta_sum_out_tmp[5][22];
        eta_sum[5][23]  = eta_sum_out_tmp[5][23];
        eta_sum[5][24]  = eta_sum_out_tmp[5][24];
        eta_sum[5][25]  = eta_sum_out_tmp[5][25];
        eta_sum[5][26]  = eta_sum_out_tmp[5][26];
        eta_sum[5][27]  = eta_sum_out_tmp[5][27];
        eta_sum[5][28]  = eta_sum_out_tmp[5][28];
        eta_sum[5][29]  = eta_sum_out_tmp[5][29];
        eta_sum[5][30]  = eta_sum_out_tmp[5][30];
        eta_sum[5][31]  = eta_sum_out_tmp[5][31];
        eta_sum[5][32]  = eta_sum_out_tmp[5][32];
        eta_sum[5][33]  = eta_sum_out_tmp[5][33];
        eta_sum[5][34]  = eta_sum_out_tmp[5][34];
        eta_sum[5][35]  = eta_sum_out_tmp[5][35];
        eta_sum[5][36]  = eta_sum_out_tmp[5][36];
        eta_sum[5][37]  = eta_sum_out_tmp[5][37];
        eta_sum[5][38]  = eta_sum_out_tmp[5][38];
        eta_sum[5][39]  = eta_sum_out_tmp[5][39];
        eta_sum[5][40]  = eta_sum_out_tmp[5][40];
        eta_sum[5][41]  = eta_sum_out_tmp[5][41];
    end
 
    1:begin 
        eta_sum[5][0]  = eta_sum_out_tmp[5][0];
        eta_sum[5][1]  = eta_sum_out_tmp[5][1];
        eta_sum[5][2]  = eta_sum_out_tmp[5][2];
        eta_sum[5][3]  = eta_sum_out_tmp[5][3];
        eta_sum[5][4]  = eta_sum_out_tmp[5][4];
        eta_sum[5][5]  = eta_sum_out_tmp[5][5];
        eta_sum[5][6]  = eta_sum_out_tmp[5][6];
        eta_sum[5][7]  = eta_sum_out_tmp[5][7];
        eta_sum[5][8]  = eta_sum_out_tmp[5][8];
        eta_sum[5][9]  = eta_sum_out_tmp[5][9];
        eta_sum[5][10]  = eta_sum_out_tmp[5][10];
        eta_sum[5][11]  = eta_sum_out_tmp[5][11];
        eta_sum[5][12]  = eta_sum_out_tmp[5][12];
        eta_sum[5][13]  = eta_sum_out_tmp[5][13];
        eta_sum[5][14]  = eta_sum_out_tmp[5][14];
        eta_sum[5][15]  = eta_sum_out_tmp[5][15];
        eta_sum[5][16]  = eta_sum_out_tmp[5][16];
        eta_sum[5][17]  = eta_sum_out_tmp[5][17];
        eta_sum[5][18]  = eta_sum_out_tmp[5][18];
        eta_sum[5][19]  = eta_sum_out_tmp[5][19];
        eta_sum[5][20]  = eta_sum_out_tmp[5][20];
        eta_sum[5][21]  = eta_sum_out_tmp[5][21];
        eta_sum[5][22]  = eta_sum_out_tmp[5][22];
        eta_sum[5][23]  = eta_sum_out_tmp[5][23];
        eta_sum[5][24]  = eta_sum_out_tmp[5][24];
        eta_sum[5][25]  = eta_sum_out_tmp[5][25];
        eta_sum[5][26]  = eta_sum_out_tmp[5][26];
        eta_sum[5][27]  = eta_sum_out_tmp[5][27];
        eta_sum[5][28]  = eta_sum_out_tmp[5][28];
        eta_sum[5][29]  = eta_sum_out_tmp[5][29];
        eta_sum[5][30]  = eta_sum_out_tmp[5][30];
        eta_sum[5][31]  = eta_sum_out_tmp[5][31];
        eta_sum[5][32]  = eta_sum_out_tmp[5][32];
        eta_sum[5][33]  = eta_sum_out_tmp[5][33];
        eta_sum[5][34]  = eta_sum_out_tmp[5][34];
        eta_sum[5][35]  = eta_sum_out_tmp[5][35];
        eta_sum[5][36]  = eta_sum_out_tmp[5][36];
        eta_sum[5][37]  = eta_sum_out_tmp[5][37];
        eta_sum[5][38]  = eta_sum_out_tmp[5][38];
        eta_sum[5][39]  = eta_sum_out_tmp[5][39];
        eta_sum[5][40]  = eta_sum_out_tmp[5][40];
        eta_sum[5][41]  = eta_sum_out_tmp[5][41];
    end
 
    2:begin 
        eta_sum[5][7]  = eta_sum_out_tmp[5][0];
        eta_sum[5][8]  = eta_sum_out_tmp[5][1];
        eta_sum[5][9]  = eta_sum_out_tmp[5][2];
        eta_sum[5][10]  = eta_sum_out_tmp[5][3];
        eta_sum[5][11]  = eta_sum_out_tmp[5][4];
        eta_sum[5][12]  = eta_sum_out_tmp[5][5];
        eta_sum[5][13]  = eta_sum_out_tmp[5][6];
        eta_sum[5][14]  = eta_sum_out_tmp[5][7];
        eta_sum[5][15]  = eta_sum_out_tmp[5][8];
        eta_sum[5][16]  = eta_sum_out_tmp[5][9];
        eta_sum[5][17]  = eta_sum_out_tmp[5][10];
        eta_sum[5][18]  = eta_sum_out_tmp[5][11];
        eta_sum[5][19]  = eta_sum_out_tmp[5][12];
        eta_sum[5][20]  = eta_sum_out_tmp[5][13];
        eta_sum[5][21]  = eta_sum_out_tmp[5][14];
        eta_sum[5][22]  = eta_sum_out_tmp[5][15];
        eta_sum[5][23]  = eta_sum_out_tmp[5][16];
        eta_sum[5][24]  = eta_sum_out_tmp[5][17];
        eta_sum[5][25]  = eta_sum_out_tmp[5][18];
        eta_sum[5][26]  = eta_sum_out_tmp[5][19];
        eta_sum[5][27]  = eta_sum_out_tmp[5][20];
        eta_sum[5][28]  = eta_sum_out_tmp[5][21];
        eta_sum[5][29]  = eta_sum_out_tmp[5][22];
        eta_sum[5][30]  = eta_sum_out_tmp[5][23];
        eta_sum[5][31]  = eta_sum_out_tmp[5][24];
        eta_sum[5][32]  = eta_sum_out_tmp[5][25];
        eta_sum[5][33]  = eta_sum_out_tmp[5][26];
        eta_sum[5][34]  = eta_sum_out_tmp[5][27];
        eta_sum[5][35]  = eta_sum_out_tmp[5][28];
        eta_sum[5][36]  = eta_sum_out_tmp[5][29];
        eta_sum[5][37]  = eta_sum_out_tmp[5][30];
        eta_sum[5][38]  = eta_sum_out_tmp[5][31];
        eta_sum[5][39]  = eta_sum_out_tmp[5][32];
        eta_sum[5][40]  = eta_sum_out_tmp[5][33];
        eta_sum[5][41]  = eta_sum_out_tmp[5][34];
        eta_sum[5][0]  = eta_sum_out_tmp[5][35];
        eta_sum[5][1]  = eta_sum_out_tmp[5][36];
        eta_sum[5][2]  = eta_sum_out_tmp[5][37];
        eta_sum[5][3]  = eta_sum_out_tmp[5][38];
        eta_sum[5][4]  = eta_sum_out_tmp[5][39];
        eta_sum[5][5]  = eta_sum_out_tmp[5][40];
        eta_sum[5][6]  = eta_sum_out_tmp[5][41];
    end
 
    3:begin 
        eta_sum[5][12]  = eta_sum_out_tmp[5][0];
        eta_sum[5][13]  = eta_sum_out_tmp[5][1];
        eta_sum[5][14]  = eta_sum_out_tmp[5][2];
        eta_sum[5][15]  = eta_sum_out_tmp[5][3];
        eta_sum[5][16]  = eta_sum_out_tmp[5][4];
        eta_sum[5][17]  = eta_sum_out_tmp[5][5];
        eta_sum[5][18]  = eta_sum_out_tmp[5][6];
        eta_sum[5][19]  = eta_sum_out_tmp[5][7];
        eta_sum[5][20]  = eta_sum_out_tmp[5][8];
        eta_sum[5][21]  = eta_sum_out_tmp[5][9];
        eta_sum[5][22]  = eta_sum_out_tmp[5][10];
        eta_sum[5][23]  = eta_sum_out_tmp[5][11];
        eta_sum[5][24]  = eta_sum_out_tmp[5][12];
        eta_sum[5][25]  = eta_sum_out_tmp[5][13];
        eta_sum[5][26]  = eta_sum_out_tmp[5][14];
        eta_sum[5][27]  = eta_sum_out_tmp[5][15];
        eta_sum[5][28]  = eta_sum_out_tmp[5][16];
        eta_sum[5][29]  = eta_sum_out_tmp[5][17];
        eta_sum[5][30]  = eta_sum_out_tmp[5][18];
        eta_sum[5][31]  = eta_sum_out_tmp[5][19];
        eta_sum[5][32]  = eta_sum_out_tmp[5][20];
        eta_sum[5][33]  = eta_sum_out_tmp[5][21];
        eta_sum[5][34]  = eta_sum_out_tmp[5][22];
        eta_sum[5][35]  = eta_sum_out_tmp[5][23];
        eta_sum[5][36]  = eta_sum_out_tmp[5][24];
        eta_sum[5][37]  = eta_sum_out_tmp[5][25];
        eta_sum[5][38]  = eta_sum_out_tmp[5][26];
        eta_sum[5][39]  = eta_sum_out_tmp[5][27];
        eta_sum[5][40]  = eta_sum_out_tmp[5][28];
        eta_sum[5][41]  = eta_sum_out_tmp[5][29];
        eta_sum[5][0]  = eta_sum_out_tmp[5][30];
        eta_sum[5][1]  = eta_sum_out_tmp[5][31];
        eta_sum[5][2]  = eta_sum_out_tmp[5][32];
        eta_sum[5][3]  = eta_sum_out_tmp[5][33];
        eta_sum[5][4]  = eta_sum_out_tmp[5][34];
        eta_sum[5][5]  = eta_sum_out_tmp[5][35];
        eta_sum[5][6]  = eta_sum_out_tmp[5][36];
        eta_sum[5][7]  = eta_sum_out_tmp[5][37];
        eta_sum[5][8]  = eta_sum_out_tmp[5][38];
        eta_sum[5][9]  = eta_sum_out_tmp[5][39];
        eta_sum[5][10]  = eta_sum_out_tmp[5][40];
        eta_sum[5][11]  = eta_sum_out_tmp[5][41];
    end
 
    4:begin 
        eta_sum[5][0]  = eta_sum_out_tmp[5][0];
        eta_sum[5][1]  = eta_sum_out_tmp[5][1];
        eta_sum[5][2]  = eta_sum_out_tmp[5][2];
        eta_sum[5][3]  = eta_sum_out_tmp[5][3];
        eta_sum[5][4]  = eta_sum_out_tmp[5][4];
        eta_sum[5][5]  = eta_sum_out_tmp[5][5];
        eta_sum[5][6]  = eta_sum_out_tmp[5][6];
        eta_sum[5][7]  = eta_sum_out_tmp[5][7];
        eta_sum[5][8]  = eta_sum_out_tmp[5][8];
        eta_sum[5][9]  = eta_sum_out_tmp[5][9];
        eta_sum[5][10]  = eta_sum_out_tmp[5][10];
        eta_sum[5][11]  = eta_sum_out_tmp[5][11];
        eta_sum[5][12]  = eta_sum_out_tmp[5][12];
        eta_sum[5][13]  = eta_sum_out_tmp[5][13];
        eta_sum[5][14]  = eta_sum_out_tmp[5][14];
        eta_sum[5][15]  = eta_sum_out_tmp[5][15];
        eta_sum[5][16]  = eta_sum_out_tmp[5][16];
        eta_sum[5][17]  = eta_sum_out_tmp[5][17];
        eta_sum[5][18]  = eta_sum_out_tmp[5][18];
        eta_sum[5][19]  = eta_sum_out_tmp[5][19];
        eta_sum[5][20]  = eta_sum_out_tmp[5][20];
        eta_sum[5][21]  = eta_sum_out_tmp[5][21];
        eta_sum[5][22]  = eta_sum_out_tmp[5][22];
        eta_sum[5][23]  = eta_sum_out_tmp[5][23];
        eta_sum[5][24]  = eta_sum_out_tmp[5][24];
        eta_sum[5][25]  = eta_sum_out_tmp[5][25];
        eta_sum[5][26]  = eta_sum_out_tmp[5][26];
        eta_sum[5][27]  = eta_sum_out_tmp[5][27];
        eta_sum[5][28]  = eta_sum_out_tmp[5][28];
        eta_sum[5][29]  = eta_sum_out_tmp[5][29];
        eta_sum[5][30]  = eta_sum_out_tmp[5][30];
        eta_sum[5][31]  = eta_sum_out_tmp[5][31];
        eta_sum[5][32]  = eta_sum_out_tmp[5][32];
        eta_sum[5][33]  = eta_sum_out_tmp[5][33];
        eta_sum[5][34]  = eta_sum_out_tmp[5][34];
        eta_sum[5][35]  = eta_sum_out_tmp[5][35];
        eta_sum[5][36]  = eta_sum_out_tmp[5][36];
        eta_sum[5][37]  = eta_sum_out_tmp[5][37];
        eta_sum[5][38]  = eta_sum_out_tmp[5][38];
        eta_sum[5][39]  = eta_sum_out_tmp[5][39];
        eta_sum[5][40]  = eta_sum_out_tmp[5][40];
        eta_sum[5][41]  = eta_sum_out_tmp[5][41];
    end
 
    5:begin 
        eta_sum[5][22]  = eta_sum_out_tmp[5][0];
        eta_sum[5][23]  = eta_sum_out_tmp[5][1];
        eta_sum[5][24]  = eta_sum_out_tmp[5][2];
        eta_sum[5][25]  = eta_sum_out_tmp[5][3];
        eta_sum[5][26]  = eta_sum_out_tmp[5][4];
        eta_sum[5][27]  = eta_sum_out_tmp[5][5];
        eta_sum[5][28]  = eta_sum_out_tmp[5][6];
        eta_sum[5][29]  = eta_sum_out_tmp[5][7];
        eta_sum[5][30]  = eta_sum_out_tmp[5][8];
        eta_sum[5][31]  = eta_sum_out_tmp[5][9];
        eta_sum[5][32]  = eta_sum_out_tmp[5][10];
        eta_sum[5][33]  = eta_sum_out_tmp[5][11];
        eta_sum[5][34]  = eta_sum_out_tmp[5][12];
        eta_sum[5][35]  = eta_sum_out_tmp[5][13];
        eta_sum[5][36]  = eta_sum_out_tmp[5][14];
        eta_sum[5][37]  = eta_sum_out_tmp[5][15];
        eta_sum[5][38]  = eta_sum_out_tmp[5][16];
        eta_sum[5][39]  = eta_sum_out_tmp[5][17];
        eta_sum[5][40]  = eta_sum_out_tmp[5][18];
        eta_sum[5][41]  = eta_sum_out_tmp[5][19];
        eta_sum[5][0]  = eta_sum_out_tmp[5][20];
        eta_sum[5][1]  = eta_sum_out_tmp[5][21];
        eta_sum[5][2]  = eta_sum_out_tmp[5][22];
        eta_sum[5][3]  = eta_sum_out_tmp[5][23];
        eta_sum[5][4]  = eta_sum_out_tmp[5][24];
        eta_sum[5][5]  = eta_sum_out_tmp[5][25];
        eta_sum[5][6]  = eta_sum_out_tmp[5][26];
        eta_sum[5][7]  = eta_sum_out_tmp[5][27];
        eta_sum[5][8]  = eta_sum_out_tmp[5][28];
        eta_sum[5][9]  = eta_sum_out_tmp[5][29];
        eta_sum[5][10]  = eta_sum_out_tmp[5][30];
        eta_sum[5][11]  = eta_sum_out_tmp[5][31];
        eta_sum[5][12]  = eta_sum_out_tmp[5][32];
        eta_sum[5][13]  = eta_sum_out_tmp[5][33];
        eta_sum[5][14]  = eta_sum_out_tmp[5][34];
        eta_sum[5][15]  = eta_sum_out_tmp[5][35];
        eta_sum[5][16]  = eta_sum_out_tmp[5][36];
        eta_sum[5][17]  = eta_sum_out_tmp[5][37];
        eta_sum[5][18]  = eta_sum_out_tmp[5][38];
        eta_sum[5][19]  = eta_sum_out_tmp[5][39];
        eta_sum[5][20]  = eta_sum_out_tmp[5][40];
        eta_sum[5][21]  = eta_sum_out_tmp[5][41];
    end
 
    6:begin 
        eta_sum[5][21]  = eta_sum_out_tmp[5][0];
        eta_sum[5][22]  = eta_sum_out_tmp[5][1];
        eta_sum[5][23]  = eta_sum_out_tmp[5][2];
        eta_sum[5][24]  = eta_sum_out_tmp[5][3];
        eta_sum[5][25]  = eta_sum_out_tmp[5][4];
        eta_sum[5][26]  = eta_sum_out_tmp[5][5];
        eta_sum[5][27]  = eta_sum_out_tmp[5][6];
        eta_sum[5][28]  = eta_sum_out_tmp[5][7];
        eta_sum[5][29]  = eta_sum_out_tmp[5][8];
        eta_sum[5][30]  = eta_sum_out_tmp[5][9];
        eta_sum[5][31]  = eta_sum_out_tmp[5][10];
        eta_sum[5][32]  = eta_sum_out_tmp[5][11];
        eta_sum[5][33]  = eta_sum_out_tmp[5][12];
        eta_sum[5][34]  = eta_sum_out_tmp[5][13];
        eta_sum[5][35]  = eta_sum_out_tmp[5][14];
        eta_sum[5][36]  = eta_sum_out_tmp[5][15];
        eta_sum[5][37]  = eta_sum_out_tmp[5][16];
        eta_sum[5][38]  = eta_sum_out_tmp[5][17];
        eta_sum[5][39]  = eta_sum_out_tmp[5][18];
        eta_sum[5][40]  = eta_sum_out_tmp[5][19];
        eta_sum[5][41]  = eta_sum_out_tmp[5][20];
        eta_sum[5][0]  = eta_sum_out_tmp[5][21];
        eta_sum[5][1]  = eta_sum_out_tmp[5][22];
        eta_sum[5][2]  = eta_sum_out_tmp[5][23];
        eta_sum[5][3]  = eta_sum_out_tmp[5][24];
        eta_sum[5][4]  = eta_sum_out_tmp[5][25];
        eta_sum[5][5]  = eta_sum_out_tmp[5][26];
        eta_sum[5][6]  = eta_sum_out_tmp[5][27];
        eta_sum[5][7]  = eta_sum_out_tmp[5][28];
        eta_sum[5][8]  = eta_sum_out_tmp[5][29];
        eta_sum[5][9]  = eta_sum_out_tmp[5][30];
        eta_sum[5][10]  = eta_sum_out_tmp[5][31];
        eta_sum[5][11]  = eta_sum_out_tmp[5][32];
        eta_sum[5][12]  = eta_sum_out_tmp[5][33];
        eta_sum[5][13]  = eta_sum_out_tmp[5][34];
        eta_sum[5][14]  = eta_sum_out_tmp[5][35];
        eta_sum[5][15]  = eta_sum_out_tmp[5][36];
        eta_sum[5][16]  = eta_sum_out_tmp[5][37];
        eta_sum[5][17]  = eta_sum_out_tmp[5][38];
        eta_sum[5][18]  = eta_sum_out_tmp[5][39];
        eta_sum[5][19]  = eta_sum_out_tmp[5][40];
        eta_sum[5][20]  = eta_sum_out_tmp[5][41];
    end
 
    7:begin 
        eta_sum[5][0]  = eta_sum_out_tmp[5][0];
        eta_sum[5][1]  = eta_sum_out_tmp[5][1];
        eta_sum[5][2]  = eta_sum_out_tmp[5][2];
        eta_sum[5][3]  = eta_sum_out_tmp[5][3];
        eta_sum[5][4]  = eta_sum_out_tmp[5][4];
        eta_sum[5][5]  = eta_sum_out_tmp[5][5];
        eta_sum[5][6]  = eta_sum_out_tmp[5][6];
        eta_sum[5][7]  = eta_sum_out_tmp[5][7];
        eta_sum[5][8]  = eta_sum_out_tmp[5][8];
        eta_sum[5][9]  = eta_sum_out_tmp[5][9];
        eta_sum[5][10]  = eta_sum_out_tmp[5][10];
        eta_sum[5][11]  = eta_sum_out_tmp[5][11];
        eta_sum[5][12]  = eta_sum_out_tmp[5][12];
        eta_sum[5][13]  = eta_sum_out_tmp[5][13];
        eta_sum[5][14]  = eta_sum_out_tmp[5][14];
        eta_sum[5][15]  = eta_sum_out_tmp[5][15];
        eta_sum[5][16]  = eta_sum_out_tmp[5][16];
        eta_sum[5][17]  = eta_sum_out_tmp[5][17];
        eta_sum[5][18]  = eta_sum_out_tmp[5][18];
        eta_sum[5][19]  = eta_sum_out_tmp[5][19];
        eta_sum[5][20]  = eta_sum_out_tmp[5][20];
        eta_sum[5][21]  = eta_sum_out_tmp[5][21];
        eta_sum[5][22]  = eta_sum_out_tmp[5][22];
        eta_sum[5][23]  = eta_sum_out_tmp[5][23];
        eta_sum[5][24]  = eta_sum_out_tmp[5][24];
        eta_sum[5][25]  = eta_sum_out_tmp[5][25];
        eta_sum[5][26]  = eta_sum_out_tmp[5][26];
        eta_sum[5][27]  = eta_sum_out_tmp[5][27];
        eta_sum[5][28]  = eta_sum_out_tmp[5][28];
        eta_sum[5][29]  = eta_sum_out_tmp[5][29];
        eta_sum[5][30]  = eta_sum_out_tmp[5][30];
        eta_sum[5][31]  = eta_sum_out_tmp[5][31];
        eta_sum[5][32]  = eta_sum_out_tmp[5][32];
        eta_sum[5][33]  = eta_sum_out_tmp[5][33];
        eta_sum[5][34]  = eta_sum_out_tmp[5][34];
        eta_sum[5][35]  = eta_sum_out_tmp[5][35];
        eta_sum[5][36]  = eta_sum_out_tmp[5][36];
        eta_sum[5][37]  = eta_sum_out_tmp[5][37];
        eta_sum[5][38]  = eta_sum_out_tmp[5][38];
        eta_sum[5][39]  = eta_sum_out_tmp[5][39];
        eta_sum[5][40]  = eta_sum_out_tmp[5][40];
        eta_sum[5][41]  = eta_sum_out_tmp[5][41];
    end
 
endcase
end

if (chk_n_output_valid[0] & active_cols[6]) begin
case (curr_layer)
    0:begin 
        eta_sum[6][5]  = eta_sum_out_tmp[6][0];
        eta_sum[6][6]  = eta_sum_out_tmp[6][1];
        eta_sum[6][7]  = eta_sum_out_tmp[6][2];
        eta_sum[6][8]  = eta_sum_out_tmp[6][3];
        eta_sum[6][9]  = eta_sum_out_tmp[6][4];
        eta_sum[6][10]  = eta_sum_out_tmp[6][5];
        eta_sum[6][11]  = eta_sum_out_tmp[6][6];
        eta_sum[6][12]  = eta_sum_out_tmp[6][7];
        eta_sum[6][13]  = eta_sum_out_tmp[6][8];
        eta_sum[6][14]  = eta_sum_out_tmp[6][9];
        eta_sum[6][15]  = eta_sum_out_tmp[6][10];
        eta_sum[6][16]  = eta_sum_out_tmp[6][11];
        eta_sum[6][17]  = eta_sum_out_tmp[6][12];
        eta_sum[6][18]  = eta_sum_out_tmp[6][13];
        eta_sum[6][19]  = eta_sum_out_tmp[6][14];
        eta_sum[6][20]  = eta_sum_out_tmp[6][15];
        eta_sum[6][21]  = eta_sum_out_tmp[6][16];
        eta_sum[6][22]  = eta_sum_out_tmp[6][17];
        eta_sum[6][23]  = eta_sum_out_tmp[6][18];
        eta_sum[6][24]  = eta_sum_out_tmp[6][19];
        eta_sum[6][25]  = eta_sum_out_tmp[6][20];
        eta_sum[6][26]  = eta_sum_out_tmp[6][21];
        eta_sum[6][27]  = eta_sum_out_tmp[6][22];
        eta_sum[6][28]  = eta_sum_out_tmp[6][23];
        eta_sum[6][29]  = eta_sum_out_tmp[6][24];
        eta_sum[6][30]  = eta_sum_out_tmp[6][25];
        eta_sum[6][31]  = eta_sum_out_tmp[6][26];
        eta_sum[6][32]  = eta_sum_out_tmp[6][27];
        eta_sum[6][33]  = eta_sum_out_tmp[6][28];
        eta_sum[6][34]  = eta_sum_out_tmp[6][29];
        eta_sum[6][35]  = eta_sum_out_tmp[6][30];
        eta_sum[6][36]  = eta_sum_out_tmp[6][31];
        eta_sum[6][37]  = eta_sum_out_tmp[6][32];
        eta_sum[6][38]  = eta_sum_out_tmp[6][33];
        eta_sum[6][39]  = eta_sum_out_tmp[6][34];
        eta_sum[6][40]  = eta_sum_out_tmp[6][35];
        eta_sum[6][41]  = eta_sum_out_tmp[6][36];
        eta_sum[6][0]  = eta_sum_out_tmp[6][37];
        eta_sum[6][1]  = eta_sum_out_tmp[6][38];
        eta_sum[6][2]  = eta_sum_out_tmp[6][39];
        eta_sum[6][3]  = eta_sum_out_tmp[6][40];
        eta_sum[6][4]  = eta_sum_out_tmp[6][41];
    end
 
    1:begin 
        eta_sum[6][0]  = eta_sum_out_tmp[6][0];
        eta_sum[6][1]  = eta_sum_out_tmp[6][1];
        eta_sum[6][2]  = eta_sum_out_tmp[6][2];
        eta_sum[6][3]  = eta_sum_out_tmp[6][3];
        eta_sum[6][4]  = eta_sum_out_tmp[6][4];
        eta_sum[6][5]  = eta_sum_out_tmp[6][5];
        eta_sum[6][6]  = eta_sum_out_tmp[6][6];
        eta_sum[6][7]  = eta_sum_out_tmp[6][7];
        eta_sum[6][8]  = eta_sum_out_tmp[6][8];
        eta_sum[6][9]  = eta_sum_out_tmp[6][9];
        eta_sum[6][10]  = eta_sum_out_tmp[6][10];
        eta_sum[6][11]  = eta_sum_out_tmp[6][11];
        eta_sum[6][12]  = eta_sum_out_tmp[6][12];
        eta_sum[6][13]  = eta_sum_out_tmp[6][13];
        eta_sum[6][14]  = eta_sum_out_tmp[6][14];
        eta_sum[6][15]  = eta_sum_out_tmp[6][15];
        eta_sum[6][16]  = eta_sum_out_tmp[6][16];
        eta_sum[6][17]  = eta_sum_out_tmp[6][17];
        eta_sum[6][18]  = eta_sum_out_tmp[6][18];
        eta_sum[6][19]  = eta_sum_out_tmp[6][19];
        eta_sum[6][20]  = eta_sum_out_tmp[6][20];
        eta_sum[6][21]  = eta_sum_out_tmp[6][21];
        eta_sum[6][22]  = eta_sum_out_tmp[6][22];
        eta_sum[6][23]  = eta_sum_out_tmp[6][23];
        eta_sum[6][24]  = eta_sum_out_tmp[6][24];
        eta_sum[6][25]  = eta_sum_out_tmp[6][25];
        eta_sum[6][26]  = eta_sum_out_tmp[6][26];
        eta_sum[6][27]  = eta_sum_out_tmp[6][27];
        eta_sum[6][28]  = eta_sum_out_tmp[6][28];
        eta_sum[6][29]  = eta_sum_out_tmp[6][29];
        eta_sum[6][30]  = eta_sum_out_tmp[6][30];
        eta_sum[6][31]  = eta_sum_out_tmp[6][31];
        eta_sum[6][32]  = eta_sum_out_tmp[6][32];
        eta_sum[6][33]  = eta_sum_out_tmp[6][33];
        eta_sum[6][34]  = eta_sum_out_tmp[6][34];
        eta_sum[6][35]  = eta_sum_out_tmp[6][35];
        eta_sum[6][36]  = eta_sum_out_tmp[6][36];
        eta_sum[6][37]  = eta_sum_out_tmp[6][37];
        eta_sum[6][38]  = eta_sum_out_tmp[6][38];
        eta_sum[6][39]  = eta_sum_out_tmp[6][39];
        eta_sum[6][40]  = eta_sum_out_tmp[6][40];
        eta_sum[6][41]  = eta_sum_out_tmp[6][41];
    end
 
    2:begin 
        eta_sum[6][0]  = eta_sum_out_tmp[6][0];
        eta_sum[6][1]  = eta_sum_out_tmp[6][1];
        eta_sum[6][2]  = eta_sum_out_tmp[6][2];
        eta_sum[6][3]  = eta_sum_out_tmp[6][3];
        eta_sum[6][4]  = eta_sum_out_tmp[6][4];
        eta_sum[6][5]  = eta_sum_out_tmp[6][5];
        eta_sum[6][6]  = eta_sum_out_tmp[6][6];
        eta_sum[6][7]  = eta_sum_out_tmp[6][7];
        eta_sum[6][8]  = eta_sum_out_tmp[6][8];
        eta_sum[6][9]  = eta_sum_out_tmp[6][9];
        eta_sum[6][10]  = eta_sum_out_tmp[6][10];
        eta_sum[6][11]  = eta_sum_out_tmp[6][11];
        eta_sum[6][12]  = eta_sum_out_tmp[6][12];
        eta_sum[6][13]  = eta_sum_out_tmp[6][13];
        eta_sum[6][14]  = eta_sum_out_tmp[6][14];
        eta_sum[6][15]  = eta_sum_out_tmp[6][15];
        eta_sum[6][16]  = eta_sum_out_tmp[6][16];
        eta_sum[6][17]  = eta_sum_out_tmp[6][17];
        eta_sum[6][18]  = eta_sum_out_tmp[6][18];
        eta_sum[6][19]  = eta_sum_out_tmp[6][19];
        eta_sum[6][20]  = eta_sum_out_tmp[6][20];
        eta_sum[6][21]  = eta_sum_out_tmp[6][21];
        eta_sum[6][22]  = eta_sum_out_tmp[6][22];
        eta_sum[6][23]  = eta_sum_out_tmp[6][23];
        eta_sum[6][24]  = eta_sum_out_tmp[6][24];
        eta_sum[6][25]  = eta_sum_out_tmp[6][25];
        eta_sum[6][26]  = eta_sum_out_tmp[6][26];
        eta_sum[6][27]  = eta_sum_out_tmp[6][27];
        eta_sum[6][28]  = eta_sum_out_tmp[6][28];
        eta_sum[6][29]  = eta_sum_out_tmp[6][29];
        eta_sum[6][30]  = eta_sum_out_tmp[6][30];
        eta_sum[6][31]  = eta_sum_out_tmp[6][31];
        eta_sum[6][32]  = eta_sum_out_tmp[6][32];
        eta_sum[6][33]  = eta_sum_out_tmp[6][33];
        eta_sum[6][34]  = eta_sum_out_tmp[6][34];
        eta_sum[6][35]  = eta_sum_out_tmp[6][35];
        eta_sum[6][36]  = eta_sum_out_tmp[6][36];
        eta_sum[6][37]  = eta_sum_out_tmp[6][37];
        eta_sum[6][38]  = eta_sum_out_tmp[6][38];
        eta_sum[6][39]  = eta_sum_out_tmp[6][39];
        eta_sum[6][40]  = eta_sum_out_tmp[6][40];
        eta_sum[6][41]  = eta_sum_out_tmp[6][41];
    end
 
    3:begin 
        eta_sum[6][20]  = eta_sum_out_tmp[6][0];
        eta_sum[6][21]  = eta_sum_out_tmp[6][1];
        eta_sum[6][22]  = eta_sum_out_tmp[6][2];
        eta_sum[6][23]  = eta_sum_out_tmp[6][3];
        eta_sum[6][24]  = eta_sum_out_tmp[6][4];
        eta_sum[6][25]  = eta_sum_out_tmp[6][5];
        eta_sum[6][26]  = eta_sum_out_tmp[6][6];
        eta_sum[6][27]  = eta_sum_out_tmp[6][7];
        eta_sum[6][28]  = eta_sum_out_tmp[6][8];
        eta_sum[6][29]  = eta_sum_out_tmp[6][9];
        eta_sum[6][30]  = eta_sum_out_tmp[6][10];
        eta_sum[6][31]  = eta_sum_out_tmp[6][11];
        eta_sum[6][32]  = eta_sum_out_tmp[6][12];
        eta_sum[6][33]  = eta_sum_out_tmp[6][13];
        eta_sum[6][34]  = eta_sum_out_tmp[6][14];
        eta_sum[6][35]  = eta_sum_out_tmp[6][15];
        eta_sum[6][36]  = eta_sum_out_tmp[6][16];
        eta_sum[6][37]  = eta_sum_out_tmp[6][17];
        eta_sum[6][38]  = eta_sum_out_tmp[6][18];
        eta_sum[6][39]  = eta_sum_out_tmp[6][19];
        eta_sum[6][40]  = eta_sum_out_tmp[6][20];
        eta_sum[6][41]  = eta_sum_out_tmp[6][21];
        eta_sum[6][0]  = eta_sum_out_tmp[6][22];
        eta_sum[6][1]  = eta_sum_out_tmp[6][23];
        eta_sum[6][2]  = eta_sum_out_tmp[6][24];
        eta_sum[6][3]  = eta_sum_out_tmp[6][25];
        eta_sum[6][4]  = eta_sum_out_tmp[6][26];
        eta_sum[6][5]  = eta_sum_out_tmp[6][27];
        eta_sum[6][6]  = eta_sum_out_tmp[6][28];
        eta_sum[6][7]  = eta_sum_out_tmp[6][29];
        eta_sum[6][8]  = eta_sum_out_tmp[6][30];
        eta_sum[6][9]  = eta_sum_out_tmp[6][31];
        eta_sum[6][10]  = eta_sum_out_tmp[6][32];
        eta_sum[6][11]  = eta_sum_out_tmp[6][33];
        eta_sum[6][12]  = eta_sum_out_tmp[6][34];
        eta_sum[6][13]  = eta_sum_out_tmp[6][35];
        eta_sum[6][14]  = eta_sum_out_tmp[6][36];
        eta_sum[6][15]  = eta_sum_out_tmp[6][37];
        eta_sum[6][16]  = eta_sum_out_tmp[6][38];
        eta_sum[6][17]  = eta_sum_out_tmp[6][39];
        eta_sum[6][18]  = eta_sum_out_tmp[6][40];
        eta_sum[6][19]  = eta_sum_out_tmp[6][41];
    end
 
    4:begin 
        eta_sum[6][39]  = eta_sum_out_tmp[6][0];
        eta_sum[6][40]  = eta_sum_out_tmp[6][1];
        eta_sum[6][41]  = eta_sum_out_tmp[6][2];
        eta_sum[6][0]  = eta_sum_out_tmp[6][3];
        eta_sum[6][1]  = eta_sum_out_tmp[6][4];
        eta_sum[6][2]  = eta_sum_out_tmp[6][5];
        eta_sum[6][3]  = eta_sum_out_tmp[6][6];
        eta_sum[6][4]  = eta_sum_out_tmp[6][7];
        eta_sum[6][5]  = eta_sum_out_tmp[6][8];
        eta_sum[6][6]  = eta_sum_out_tmp[6][9];
        eta_sum[6][7]  = eta_sum_out_tmp[6][10];
        eta_sum[6][8]  = eta_sum_out_tmp[6][11];
        eta_sum[6][9]  = eta_sum_out_tmp[6][12];
        eta_sum[6][10]  = eta_sum_out_tmp[6][13];
        eta_sum[6][11]  = eta_sum_out_tmp[6][14];
        eta_sum[6][12]  = eta_sum_out_tmp[6][15];
        eta_sum[6][13]  = eta_sum_out_tmp[6][16];
        eta_sum[6][14]  = eta_sum_out_tmp[6][17];
        eta_sum[6][15]  = eta_sum_out_tmp[6][18];
        eta_sum[6][16]  = eta_sum_out_tmp[6][19];
        eta_sum[6][17]  = eta_sum_out_tmp[6][20];
        eta_sum[6][18]  = eta_sum_out_tmp[6][21];
        eta_sum[6][19]  = eta_sum_out_tmp[6][22];
        eta_sum[6][20]  = eta_sum_out_tmp[6][23];
        eta_sum[6][21]  = eta_sum_out_tmp[6][24];
        eta_sum[6][22]  = eta_sum_out_tmp[6][25];
        eta_sum[6][23]  = eta_sum_out_tmp[6][26];
        eta_sum[6][24]  = eta_sum_out_tmp[6][27];
        eta_sum[6][25]  = eta_sum_out_tmp[6][28];
        eta_sum[6][26]  = eta_sum_out_tmp[6][29];
        eta_sum[6][27]  = eta_sum_out_tmp[6][30];
        eta_sum[6][28]  = eta_sum_out_tmp[6][31];
        eta_sum[6][29]  = eta_sum_out_tmp[6][32];
        eta_sum[6][30]  = eta_sum_out_tmp[6][33];
        eta_sum[6][31]  = eta_sum_out_tmp[6][34];
        eta_sum[6][32]  = eta_sum_out_tmp[6][35];
        eta_sum[6][33]  = eta_sum_out_tmp[6][36];
        eta_sum[6][34]  = eta_sum_out_tmp[6][37];
        eta_sum[6][35]  = eta_sum_out_tmp[6][38];
        eta_sum[6][36]  = eta_sum_out_tmp[6][39];
        eta_sum[6][37]  = eta_sum_out_tmp[6][40];
        eta_sum[6][38]  = eta_sum_out_tmp[6][41];
    end
 
    5:begin 
        eta_sum[6][0]  = eta_sum_out_tmp[6][0];
        eta_sum[6][1]  = eta_sum_out_tmp[6][1];
        eta_sum[6][2]  = eta_sum_out_tmp[6][2];
        eta_sum[6][3]  = eta_sum_out_tmp[6][3];
        eta_sum[6][4]  = eta_sum_out_tmp[6][4];
        eta_sum[6][5]  = eta_sum_out_tmp[6][5];
        eta_sum[6][6]  = eta_sum_out_tmp[6][6];
        eta_sum[6][7]  = eta_sum_out_tmp[6][7];
        eta_sum[6][8]  = eta_sum_out_tmp[6][8];
        eta_sum[6][9]  = eta_sum_out_tmp[6][9];
        eta_sum[6][10]  = eta_sum_out_tmp[6][10];
        eta_sum[6][11]  = eta_sum_out_tmp[6][11];
        eta_sum[6][12]  = eta_sum_out_tmp[6][12];
        eta_sum[6][13]  = eta_sum_out_tmp[6][13];
        eta_sum[6][14]  = eta_sum_out_tmp[6][14];
        eta_sum[6][15]  = eta_sum_out_tmp[6][15];
        eta_sum[6][16]  = eta_sum_out_tmp[6][16];
        eta_sum[6][17]  = eta_sum_out_tmp[6][17];
        eta_sum[6][18]  = eta_sum_out_tmp[6][18];
        eta_sum[6][19]  = eta_sum_out_tmp[6][19];
        eta_sum[6][20]  = eta_sum_out_tmp[6][20];
        eta_sum[6][21]  = eta_sum_out_tmp[6][21];
        eta_sum[6][22]  = eta_sum_out_tmp[6][22];
        eta_sum[6][23]  = eta_sum_out_tmp[6][23];
        eta_sum[6][24]  = eta_sum_out_tmp[6][24];
        eta_sum[6][25]  = eta_sum_out_tmp[6][25];
        eta_sum[6][26]  = eta_sum_out_tmp[6][26];
        eta_sum[6][27]  = eta_sum_out_tmp[6][27];
        eta_sum[6][28]  = eta_sum_out_tmp[6][28];
        eta_sum[6][29]  = eta_sum_out_tmp[6][29];
        eta_sum[6][30]  = eta_sum_out_tmp[6][30];
        eta_sum[6][31]  = eta_sum_out_tmp[6][31];
        eta_sum[6][32]  = eta_sum_out_tmp[6][32];
        eta_sum[6][33]  = eta_sum_out_tmp[6][33];
        eta_sum[6][34]  = eta_sum_out_tmp[6][34];
        eta_sum[6][35]  = eta_sum_out_tmp[6][35];
        eta_sum[6][36]  = eta_sum_out_tmp[6][36];
        eta_sum[6][37]  = eta_sum_out_tmp[6][37];
        eta_sum[6][38]  = eta_sum_out_tmp[6][38];
        eta_sum[6][39]  = eta_sum_out_tmp[6][39];
        eta_sum[6][40]  = eta_sum_out_tmp[6][40];
        eta_sum[6][41]  = eta_sum_out_tmp[6][41];
    end
 
    6:begin 
        eta_sum[6][0]  = eta_sum_out_tmp[6][0];
        eta_sum[6][1]  = eta_sum_out_tmp[6][1];
        eta_sum[6][2]  = eta_sum_out_tmp[6][2];
        eta_sum[6][3]  = eta_sum_out_tmp[6][3];
        eta_sum[6][4]  = eta_sum_out_tmp[6][4];
        eta_sum[6][5]  = eta_sum_out_tmp[6][5];
        eta_sum[6][6]  = eta_sum_out_tmp[6][6];
        eta_sum[6][7]  = eta_sum_out_tmp[6][7];
        eta_sum[6][8]  = eta_sum_out_tmp[6][8];
        eta_sum[6][9]  = eta_sum_out_tmp[6][9];
        eta_sum[6][10]  = eta_sum_out_tmp[6][10];
        eta_sum[6][11]  = eta_sum_out_tmp[6][11];
        eta_sum[6][12]  = eta_sum_out_tmp[6][12];
        eta_sum[6][13]  = eta_sum_out_tmp[6][13];
        eta_sum[6][14]  = eta_sum_out_tmp[6][14];
        eta_sum[6][15]  = eta_sum_out_tmp[6][15];
        eta_sum[6][16]  = eta_sum_out_tmp[6][16];
        eta_sum[6][17]  = eta_sum_out_tmp[6][17];
        eta_sum[6][18]  = eta_sum_out_tmp[6][18];
        eta_sum[6][19]  = eta_sum_out_tmp[6][19];
        eta_sum[6][20]  = eta_sum_out_tmp[6][20];
        eta_sum[6][21]  = eta_sum_out_tmp[6][21];
        eta_sum[6][22]  = eta_sum_out_tmp[6][22];
        eta_sum[6][23]  = eta_sum_out_tmp[6][23];
        eta_sum[6][24]  = eta_sum_out_tmp[6][24];
        eta_sum[6][25]  = eta_sum_out_tmp[6][25];
        eta_sum[6][26]  = eta_sum_out_tmp[6][26];
        eta_sum[6][27]  = eta_sum_out_tmp[6][27];
        eta_sum[6][28]  = eta_sum_out_tmp[6][28];
        eta_sum[6][29]  = eta_sum_out_tmp[6][29];
        eta_sum[6][30]  = eta_sum_out_tmp[6][30];
        eta_sum[6][31]  = eta_sum_out_tmp[6][31];
        eta_sum[6][32]  = eta_sum_out_tmp[6][32];
        eta_sum[6][33]  = eta_sum_out_tmp[6][33];
        eta_sum[6][34]  = eta_sum_out_tmp[6][34];
        eta_sum[6][35]  = eta_sum_out_tmp[6][35];
        eta_sum[6][36]  = eta_sum_out_tmp[6][36];
        eta_sum[6][37]  = eta_sum_out_tmp[6][37];
        eta_sum[6][38]  = eta_sum_out_tmp[6][38];
        eta_sum[6][39]  = eta_sum_out_tmp[6][39];
        eta_sum[6][40]  = eta_sum_out_tmp[6][40];
        eta_sum[6][41]  = eta_sum_out_tmp[6][41];
    end
 
    7:begin 
        eta_sum[6][14]  = eta_sum_out_tmp[6][0];
        eta_sum[6][15]  = eta_sum_out_tmp[6][1];
        eta_sum[6][16]  = eta_sum_out_tmp[6][2];
        eta_sum[6][17]  = eta_sum_out_tmp[6][3];
        eta_sum[6][18]  = eta_sum_out_tmp[6][4];
        eta_sum[6][19]  = eta_sum_out_tmp[6][5];
        eta_sum[6][20]  = eta_sum_out_tmp[6][6];
        eta_sum[6][21]  = eta_sum_out_tmp[6][7];
        eta_sum[6][22]  = eta_sum_out_tmp[6][8];
        eta_sum[6][23]  = eta_sum_out_tmp[6][9];
        eta_sum[6][24]  = eta_sum_out_tmp[6][10];
        eta_sum[6][25]  = eta_sum_out_tmp[6][11];
        eta_sum[6][26]  = eta_sum_out_tmp[6][12];
        eta_sum[6][27]  = eta_sum_out_tmp[6][13];
        eta_sum[6][28]  = eta_sum_out_tmp[6][14];
        eta_sum[6][29]  = eta_sum_out_tmp[6][15];
        eta_sum[6][30]  = eta_sum_out_tmp[6][16];
        eta_sum[6][31]  = eta_sum_out_tmp[6][17];
        eta_sum[6][32]  = eta_sum_out_tmp[6][18];
        eta_sum[6][33]  = eta_sum_out_tmp[6][19];
        eta_sum[6][34]  = eta_sum_out_tmp[6][20];
        eta_sum[6][35]  = eta_sum_out_tmp[6][21];
        eta_sum[6][36]  = eta_sum_out_tmp[6][22];
        eta_sum[6][37]  = eta_sum_out_tmp[6][23];
        eta_sum[6][38]  = eta_sum_out_tmp[6][24];
        eta_sum[6][39]  = eta_sum_out_tmp[6][25];
        eta_sum[6][40]  = eta_sum_out_tmp[6][26];
        eta_sum[6][41]  = eta_sum_out_tmp[6][27];
        eta_sum[6][0]  = eta_sum_out_tmp[6][28];
        eta_sum[6][1]  = eta_sum_out_tmp[6][29];
        eta_sum[6][2]  = eta_sum_out_tmp[6][30];
        eta_sum[6][3]  = eta_sum_out_tmp[6][31];
        eta_sum[6][4]  = eta_sum_out_tmp[6][32];
        eta_sum[6][5]  = eta_sum_out_tmp[6][33];
        eta_sum[6][6]  = eta_sum_out_tmp[6][34];
        eta_sum[6][7]  = eta_sum_out_tmp[6][35];
        eta_sum[6][8]  = eta_sum_out_tmp[6][36];
        eta_sum[6][9]  = eta_sum_out_tmp[6][37];
        eta_sum[6][10]  = eta_sum_out_tmp[6][38];
        eta_sum[6][11]  = eta_sum_out_tmp[6][39];
        eta_sum[6][12]  = eta_sum_out_tmp[6][40];
        eta_sum[6][13]  = eta_sum_out_tmp[6][41];
    end
 
endcase
end

if (chk_n_output_valid[0] & active_cols[7]) begin
case (curr_layer)
    0:begin 
        eta_sum[7][0]  = eta_sum_out_tmp[7][0];
        eta_sum[7][1]  = eta_sum_out_tmp[7][1];
        eta_sum[7][2]  = eta_sum_out_tmp[7][2];
        eta_sum[7][3]  = eta_sum_out_tmp[7][3];
        eta_sum[7][4]  = eta_sum_out_tmp[7][4];
        eta_sum[7][5]  = eta_sum_out_tmp[7][5];
        eta_sum[7][6]  = eta_sum_out_tmp[7][6];
        eta_sum[7][7]  = eta_sum_out_tmp[7][7];
        eta_sum[7][8]  = eta_sum_out_tmp[7][8];
        eta_sum[7][9]  = eta_sum_out_tmp[7][9];
        eta_sum[7][10]  = eta_sum_out_tmp[7][10];
        eta_sum[7][11]  = eta_sum_out_tmp[7][11];
        eta_sum[7][12]  = eta_sum_out_tmp[7][12];
        eta_sum[7][13]  = eta_sum_out_tmp[7][13];
        eta_sum[7][14]  = eta_sum_out_tmp[7][14];
        eta_sum[7][15]  = eta_sum_out_tmp[7][15];
        eta_sum[7][16]  = eta_sum_out_tmp[7][16];
        eta_sum[7][17]  = eta_sum_out_tmp[7][17];
        eta_sum[7][18]  = eta_sum_out_tmp[7][18];
        eta_sum[7][19]  = eta_sum_out_tmp[7][19];
        eta_sum[7][20]  = eta_sum_out_tmp[7][20];
        eta_sum[7][21]  = eta_sum_out_tmp[7][21];
        eta_sum[7][22]  = eta_sum_out_tmp[7][22];
        eta_sum[7][23]  = eta_sum_out_tmp[7][23];
        eta_sum[7][24]  = eta_sum_out_tmp[7][24];
        eta_sum[7][25]  = eta_sum_out_tmp[7][25];
        eta_sum[7][26]  = eta_sum_out_tmp[7][26];
        eta_sum[7][27]  = eta_sum_out_tmp[7][27];
        eta_sum[7][28]  = eta_sum_out_tmp[7][28];
        eta_sum[7][29]  = eta_sum_out_tmp[7][29];
        eta_sum[7][30]  = eta_sum_out_tmp[7][30];
        eta_sum[7][31]  = eta_sum_out_tmp[7][31];
        eta_sum[7][32]  = eta_sum_out_tmp[7][32];
        eta_sum[7][33]  = eta_sum_out_tmp[7][33];
        eta_sum[7][34]  = eta_sum_out_tmp[7][34];
        eta_sum[7][35]  = eta_sum_out_tmp[7][35];
        eta_sum[7][36]  = eta_sum_out_tmp[7][36];
        eta_sum[7][37]  = eta_sum_out_tmp[7][37];
        eta_sum[7][38]  = eta_sum_out_tmp[7][38];
        eta_sum[7][39]  = eta_sum_out_tmp[7][39];
        eta_sum[7][40]  = eta_sum_out_tmp[7][40];
        eta_sum[7][41]  = eta_sum_out_tmp[7][41];
    end
 
    1:begin 
        eta_sum[7][30]  = eta_sum_out_tmp[7][0];
        eta_sum[7][31]  = eta_sum_out_tmp[7][1];
        eta_sum[7][32]  = eta_sum_out_tmp[7][2];
        eta_sum[7][33]  = eta_sum_out_tmp[7][3];
        eta_sum[7][34]  = eta_sum_out_tmp[7][4];
        eta_sum[7][35]  = eta_sum_out_tmp[7][5];
        eta_sum[7][36]  = eta_sum_out_tmp[7][6];
        eta_sum[7][37]  = eta_sum_out_tmp[7][7];
        eta_sum[7][38]  = eta_sum_out_tmp[7][8];
        eta_sum[7][39]  = eta_sum_out_tmp[7][9];
        eta_sum[7][40]  = eta_sum_out_tmp[7][10];
        eta_sum[7][41]  = eta_sum_out_tmp[7][11];
        eta_sum[7][0]  = eta_sum_out_tmp[7][12];
        eta_sum[7][1]  = eta_sum_out_tmp[7][13];
        eta_sum[7][2]  = eta_sum_out_tmp[7][14];
        eta_sum[7][3]  = eta_sum_out_tmp[7][15];
        eta_sum[7][4]  = eta_sum_out_tmp[7][16];
        eta_sum[7][5]  = eta_sum_out_tmp[7][17];
        eta_sum[7][6]  = eta_sum_out_tmp[7][18];
        eta_sum[7][7]  = eta_sum_out_tmp[7][19];
        eta_sum[7][8]  = eta_sum_out_tmp[7][20];
        eta_sum[7][9]  = eta_sum_out_tmp[7][21];
        eta_sum[7][10]  = eta_sum_out_tmp[7][22];
        eta_sum[7][11]  = eta_sum_out_tmp[7][23];
        eta_sum[7][12]  = eta_sum_out_tmp[7][24];
        eta_sum[7][13]  = eta_sum_out_tmp[7][25];
        eta_sum[7][14]  = eta_sum_out_tmp[7][26];
        eta_sum[7][15]  = eta_sum_out_tmp[7][27];
        eta_sum[7][16]  = eta_sum_out_tmp[7][28];
        eta_sum[7][17]  = eta_sum_out_tmp[7][29];
        eta_sum[7][18]  = eta_sum_out_tmp[7][30];
        eta_sum[7][19]  = eta_sum_out_tmp[7][31];
        eta_sum[7][20]  = eta_sum_out_tmp[7][32];
        eta_sum[7][21]  = eta_sum_out_tmp[7][33];
        eta_sum[7][22]  = eta_sum_out_tmp[7][34];
        eta_sum[7][23]  = eta_sum_out_tmp[7][35];
        eta_sum[7][24]  = eta_sum_out_tmp[7][36];
        eta_sum[7][25]  = eta_sum_out_tmp[7][37];
        eta_sum[7][26]  = eta_sum_out_tmp[7][38];
        eta_sum[7][27]  = eta_sum_out_tmp[7][39];
        eta_sum[7][28]  = eta_sum_out_tmp[7][40];
        eta_sum[7][29]  = eta_sum_out_tmp[7][41];
    end
 
    2:begin 
        eta_sum[7][34]  = eta_sum_out_tmp[7][0];
        eta_sum[7][35]  = eta_sum_out_tmp[7][1];
        eta_sum[7][36]  = eta_sum_out_tmp[7][2];
        eta_sum[7][37]  = eta_sum_out_tmp[7][3];
        eta_sum[7][38]  = eta_sum_out_tmp[7][4];
        eta_sum[7][39]  = eta_sum_out_tmp[7][5];
        eta_sum[7][40]  = eta_sum_out_tmp[7][6];
        eta_sum[7][41]  = eta_sum_out_tmp[7][7];
        eta_sum[7][0]  = eta_sum_out_tmp[7][8];
        eta_sum[7][1]  = eta_sum_out_tmp[7][9];
        eta_sum[7][2]  = eta_sum_out_tmp[7][10];
        eta_sum[7][3]  = eta_sum_out_tmp[7][11];
        eta_sum[7][4]  = eta_sum_out_tmp[7][12];
        eta_sum[7][5]  = eta_sum_out_tmp[7][13];
        eta_sum[7][6]  = eta_sum_out_tmp[7][14];
        eta_sum[7][7]  = eta_sum_out_tmp[7][15];
        eta_sum[7][8]  = eta_sum_out_tmp[7][16];
        eta_sum[7][9]  = eta_sum_out_tmp[7][17];
        eta_sum[7][10]  = eta_sum_out_tmp[7][18];
        eta_sum[7][11]  = eta_sum_out_tmp[7][19];
        eta_sum[7][12]  = eta_sum_out_tmp[7][20];
        eta_sum[7][13]  = eta_sum_out_tmp[7][21];
        eta_sum[7][14]  = eta_sum_out_tmp[7][22];
        eta_sum[7][15]  = eta_sum_out_tmp[7][23];
        eta_sum[7][16]  = eta_sum_out_tmp[7][24];
        eta_sum[7][17]  = eta_sum_out_tmp[7][25];
        eta_sum[7][18]  = eta_sum_out_tmp[7][26];
        eta_sum[7][19]  = eta_sum_out_tmp[7][27];
        eta_sum[7][20]  = eta_sum_out_tmp[7][28];
        eta_sum[7][21]  = eta_sum_out_tmp[7][29];
        eta_sum[7][22]  = eta_sum_out_tmp[7][30];
        eta_sum[7][23]  = eta_sum_out_tmp[7][31];
        eta_sum[7][24]  = eta_sum_out_tmp[7][32];
        eta_sum[7][25]  = eta_sum_out_tmp[7][33];
        eta_sum[7][26]  = eta_sum_out_tmp[7][34];
        eta_sum[7][27]  = eta_sum_out_tmp[7][35];
        eta_sum[7][28]  = eta_sum_out_tmp[7][36];
        eta_sum[7][29]  = eta_sum_out_tmp[7][37];
        eta_sum[7][30]  = eta_sum_out_tmp[7][38];
        eta_sum[7][31]  = eta_sum_out_tmp[7][39];
        eta_sum[7][32]  = eta_sum_out_tmp[7][40];
        eta_sum[7][33]  = eta_sum_out_tmp[7][41];
    end
 
    3:begin 
        eta_sum[7][0]  = eta_sum_out_tmp[7][0];
        eta_sum[7][1]  = eta_sum_out_tmp[7][1];
        eta_sum[7][2]  = eta_sum_out_tmp[7][2];
        eta_sum[7][3]  = eta_sum_out_tmp[7][3];
        eta_sum[7][4]  = eta_sum_out_tmp[7][4];
        eta_sum[7][5]  = eta_sum_out_tmp[7][5];
        eta_sum[7][6]  = eta_sum_out_tmp[7][6];
        eta_sum[7][7]  = eta_sum_out_tmp[7][7];
        eta_sum[7][8]  = eta_sum_out_tmp[7][8];
        eta_sum[7][9]  = eta_sum_out_tmp[7][9];
        eta_sum[7][10]  = eta_sum_out_tmp[7][10];
        eta_sum[7][11]  = eta_sum_out_tmp[7][11];
        eta_sum[7][12]  = eta_sum_out_tmp[7][12];
        eta_sum[7][13]  = eta_sum_out_tmp[7][13];
        eta_sum[7][14]  = eta_sum_out_tmp[7][14];
        eta_sum[7][15]  = eta_sum_out_tmp[7][15];
        eta_sum[7][16]  = eta_sum_out_tmp[7][16];
        eta_sum[7][17]  = eta_sum_out_tmp[7][17];
        eta_sum[7][18]  = eta_sum_out_tmp[7][18];
        eta_sum[7][19]  = eta_sum_out_tmp[7][19];
        eta_sum[7][20]  = eta_sum_out_tmp[7][20];
        eta_sum[7][21]  = eta_sum_out_tmp[7][21];
        eta_sum[7][22]  = eta_sum_out_tmp[7][22];
        eta_sum[7][23]  = eta_sum_out_tmp[7][23];
        eta_sum[7][24]  = eta_sum_out_tmp[7][24];
        eta_sum[7][25]  = eta_sum_out_tmp[7][25];
        eta_sum[7][26]  = eta_sum_out_tmp[7][26];
        eta_sum[7][27]  = eta_sum_out_tmp[7][27];
        eta_sum[7][28]  = eta_sum_out_tmp[7][28];
        eta_sum[7][29]  = eta_sum_out_tmp[7][29];
        eta_sum[7][30]  = eta_sum_out_tmp[7][30];
        eta_sum[7][31]  = eta_sum_out_tmp[7][31];
        eta_sum[7][32]  = eta_sum_out_tmp[7][32];
        eta_sum[7][33]  = eta_sum_out_tmp[7][33];
        eta_sum[7][34]  = eta_sum_out_tmp[7][34];
        eta_sum[7][35]  = eta_sum_out_tmp[7][35];
        eta_sum[7][36]  = eta_sum_out_tmp[7][36];
        eta_sum[7][37]  = eta_sum_out_tmp[7][37];
        eta_sum[7][38]  = eta_sum_out_tmp[7][38];
        eta_sum[7][39]  = eta_sum_out_tmp[7][39];
        eta_sum[7][40]  = eta_sum_out_tmp[7][40];
        eta_sum[7][41]  = eta_sum_out_tmp[7][41];
    end
 
    4:begin 
        eta_sum[7][0]  = eta_sum_out_tmp[7][0];
        eta_sum[7][1]  = eta_sum_out_tmp[7][1];
        eta_sum[7][2]  = eta_sum_out_tmp[7][2];
        eta_sum[7][3]  = eta_sum_out_tmp[7][3];
        eta_sum[7][4]  = eta_sum_out_tmp[7][4];
        eta_sum[7][5]  = eta_sum_out_tmp[7][5];
        eta_sum[7][6]  = eta_sum_out_tmp[7][6];
        eta_sum[7][7]  = eta_sum_out_tmp[7][7];
        eta_sum[7][8]  = eta_sum_out_tmp[7][8];
        eta_sum[7][9]  = eta_sum_out_tmp[7][9];
        eta_sum[7][10]  = eta_sum_out_tmp[7][10];
        eta_sum[7][11]  = eta_sum_out_tmp[7][11];
        eta_sum[7][12]  = eta_sum_out_tmp[7][12];
        eta_sum[7][13]  = eta_sum_out_tmp[7][13];
        eta_sum[7][14]  = eta_sum_out_tmp[7][14];
        eta_sum[7][15]  = eta_sum_out_tmp[7][15];
        eta_sum[7][16]  = eta_sum_out_tmp[7][16];
        eta_sum[7][17]  = eta_sum_out_tmp[7][17];
        eta_sum[7][18]  = eta_sum_out_tmp[7][18];
        eta_sum[7][19]  = eta_sum_out_tmp[7][19];
        eta_sum[7][20]  = eta_sum_out_tmp[7][20];
        eta_sum[7][21]  = eta_sum_out_tmp[7][21];
        eta_sum[7][22]  = eta_sum_out_tmp[7][22];
        eta_sum[7][23]  = eta_sum_out_tmp[7][23];
        eta_sum[7][24]  = eta_sum_out_tmp[7][24];
        eta_sum[7][25]  = eta_sum_out_tmp[7][25];
        eta_sum[7][26]  = eta_sum_out_tmp[7][26];
        eta_sum[7][27]  = eta_sum_out_tmp[7][27];
        eta_sum[7][28]  = eta_sum_out_tmp[7][28];
        eta_sum[7][29]  = eta_sum_out_tmp[7][29];
        eta_sum[7][30]  = eta_sum_out_tmp[7][30];
        eta_sum[7][31]  = eta_sum_out_tmp[7][31];
        eta_sum[7][32]  = eta_sum_out_tmp[7][32];
        eta_sum[7][33]  = eta_sum_out_tmp[7][33];
        eta_sum[7][34]  = eta_sum_out_tmp[7][34];
        eta_sum[7][35]  = eta_sum_out_tmp[7][35];
        eta_sum[7][36]  = eta_sum_out_tmp[7][36];
        eta_sum[7][37]  = eta_sum_out_tmp[7][37];
        eta_sum[7][38]  = eta_sum_out_tmp[7][38];
        eta_sum[7][39]  = eta_sum_out_tmp[7][39];
        eta_sum[7][40]  = eta_sum_out_tmp[7][40];
        eta_sum[7][41]  = eta_sum_out_tmp[7][41];
    end
 
    5:begin 
        eta_sum[7][4]  = eta_sum_out_tmp[7][0];
        eta_sum[7][5]  = eta_sum_out_tmp[7][1];
        eta_sum[7][6]  = eta_sum_out_tmp[7][2];
        eta_sum[7][7]  = eta_sum_out_tmp[7][3];
        eta_sum[7][8]  = eta_sum_out_tmp[7][4];
        eta_sum[7][9]  = eta_sum_out_tmp[7][5];
        eta_sum[7][10]  = eta_sum_out_tmp[7][6];
        eta_sum[7][11]  = eta_sum_out_tmp[7][7];
        eta_sum[7][12]  = eta_sum_out_tmp[7][8];
        eta_sum[7][13]  = eta_sum_out_tmp[7][9];
        eta_sum[7][14]  = eta_sum_out_tmp[7][10];
        eta_sum[7][15]  = eta_sum_out_tmp[7][11];
        eta_sum[7][16]  = eta_sum_out_tmp[7][12];
        eta_sum[7][17]  = eta_sum_out_tmp[7][13];
        eta_sum[7][18]  = eta_sum_out_tmp[7][14];
        eta_sum[7][19]  = eta_sum_out_tmp[7][15];
        eta_sum[7][20]  = eta_sum_out_tmp[7][16];
        eta_sum[7][21]  = eta_sum_out_tmp[7][17];
        eta_sum[7][22]  = eta_sum_out_tmp[7][18];
        eta_sum[7][23]  = eta_sum_out_tmp[7][19];
        eta_sum[7][24]  = eta_sum_out_tmp[7][20];
        eta_sum[7][25]  = eta_sum_out_tmp[7][21];
        eta_sum[7][26]  = eta_sum_out_tmp[7][22];
        eta_sum[7][27]  = eta_sum_out_tmp[7][23];
        eta_sum[7][28]  = eta_sum_out_tmp[7][24];
        eta_sum[7][29]  = eta_sum_out_tmp[7][25];
        eta_sum[7][30]  = eta_sum_out_tmp[7][26];
        eta_sum[7][31]  = eta_sum_out_tmp[7][27];
        eta_sum[7][32]  = eta_sum_out_tmp[7][28];
        eta_sum[7][33]  = eta_sum_out_tmp[7][29];
        eta_sum[7][34]  = eta_sum_out_tmp[7][30];
        eta_sum[7][35]  = eta_sum_out_tmp[7][31];
        eta_sum[7][36]  = eta_sum_out_tmp[7][32];
        eta_sum[7][37]  = eta_sum_out_tmp[7][33];
        eta_sum[7][38]  = eta_sum_out_tmp[7][34];
        eta_sum[7][39]  = eta_sum_out_tmp[7][35];
        eta_sum[7][40]  = eta_sum_out_tmp[7][36];
        eta_sum[7][41]  = eta_sum_out_tmp[7][37];
        eta_sum[7][0]  = eta_sum_out_tmp[7][38];
        eta_sum[7][1]  = eta_sum_out_tmp[7][39];
        eta_sum[7][2]  = eta_sum_out_tmp[7][40];
        eta_sum[7][3]  = eta_sum_out_tmp[7][41];
    end
 
    6:begin 
        eta_sum[7][20]  = eta_sum_out_tmp[7][0];
        eta_sum[7][21]  = eta_sum_out_tmp[7][1];
        eta_sum[7][22]  = eta_sum_out_tmp[7][2];
        eta_sum[7][23]  = eta_sum_out_tmp[7][3];
        eta_sum[7][24]  = eta_sum_out_tmp[7][4];
        eta_sum[7][25]  = eta_sum_out_tmp[7][5];
        eta_sum[7][26]  = eta_sum_out_tmp[7][6];
        eta_sum[7][27]  = eta_sum_out_tmp[7][7];
        eta_sum[7][28]  = eta_sum_out_tmp[7][8];
        eta_sum[7][29]  = eta_sum_out_tmp[7][9];
        eta_sum[7][30]  = eta_sum_out_tmp[7][10];
        eta_sum[7][31]  = eta_sum_out_tmp[7][11];
        eta_sum[7][32]  = eta_sum_out_tmp[7][12];
        eta_sum[7][33]  = eta_sum_out_tmp[7][13];
        eta_sum[7][34]  = eta_sum_out_tmp[7][14];
        eta_sum[7][35]  = eta_sum_out_tmp[7][15];
        eta_sum[7][36]  = eta_sum_out_tmp[7][16];
        eta_sum[7][37]  = eta_sum_out_tmp[7][17];
        eta_sum[7][38]  = eta_sum_out_tmp[7][18];
        eta_sum[7][39]  = eta_sum_out_tmp[7][19];
        eta_sum[7][40]  = eta_sum_out_tmp[7][20];
        eta_sum[7][41]  = eta_sum_out_tmp[7][21];
        eta_sum[7][0]  = eta_sum_out_tmp[7][22];
        eta_sum[7][1]  = eta_sum_out_tmp[7][23];
        eta_sum[7][2]  = eta_sum_out_tmp[7][24];
        eta_sum[7][3]  = eta_sum_out_tmp[7][25];
        eta_sum[7][4]  = eta_sum_out_tmp[7][26];
        eta_sum[7][5]  = eta_sum_out_tmp[7][27];
        eta_sum[7][6]  = eta_sum_out_tmp[7][28];
        eta_sum[7][7]  = eta_sum_out_tmp[7][29];
        eta_sum[7][8]  = eta_sum_out_tmp[7][30];
        eta_sum[7][9]  = eta_sum_out_tmp[7][31];
        eta_sum[7][10]  = eta_sum_out_tmp[7][32];
        eta_sum[7][11]  = eta_sum_out_tmp[7][33];
        eta_sum[7][12]  = eta_sum_out_tmp[7][34];
        eta_sum[7][13]  = eta_sum_out_tmp[7][35];
        eta_sum[7][14]  = eta_sum_out_tmp[7][36];
        eta_sum[7][15]  = eta_sum_out_tmp[7][37];
        eta_sum[7][16]  = eta_sum_out_tmp[7][38];
        eta_sum[7][17]  = eta_sum_out_tmp[7][39];
        eta_sum[7][18]  = eta_sum_out_tmp[7][40];
        eta_sum[7][19]  = eta_sum_out_tmp[7][41];
    end
 
    7:begin 
        eta_sum[7][0]  = eta_sum_out_tmp[7][0];
        eta_sum[7][1]  = eta_sum_out_tmp[7][1];
        eta_sum[7][2]  = eta_sum_out_tmp[7][2];
        eta_sum[7][3]  = eta_sum_out_tmp[7][3];
        eta_sum[7][4]  = eta_sum_out_tmp[7][4];
        eta_sum[7][5]  = eta_sum_out_tmp[7][5];
        eta_sum[7][6]  = eta_sum_out_tmp[7][6];
        eta_sum[7][7]  = eta_sum_out_tmp[7][7];
        eta_sum[7][8]  = eta_sum_out_tmp[7][8];
        eta_sum[7][9]  = eta_sum_out_tmp[7][9];
        eta_sum[7][10]  = eta_sum_out_tmp[7][10];
        eta_sum[7][11]  = eta_sum_out_tmp[7][11];
        eta_sum[7][12]  = eta_sum_out_tmp[7][12];
        eta_sum[7][13]  = eta_sum_out_tmp[7][13];
        eta_sum[7][14]  = eta_sum_out_tmp[7][14];
        eta_sum[7][15]  = eta_sum_out_tmp[7][15];
        eta_sum[7][16]  = eta_sum_out_tmp[7][16];
        eta_sum[7][17]  = eta_sum_out_tmp[7][17];
        eta_sum[7][18]  = eta_sum_out_tmp[7][18];
        eta_sum[7][19]  = eta_sum_out_tmp[7][19];
        eta_sum[7][20]  = eta_sum_out_tmp[7][20];
        eta_sum[7][21]  = eta_sum_out_tmp[7][21];
        eta_sum[7][22]  = eta_sum_out_tmp[7][22];
        eta_sum[7][23]  = eta_sum_out_tmp[7][23];
        eta_sum[7][24]  = eta_sum_out_tmp[7][24];
        eta_sum[7][25]  = eta_sum_out_tmp[7][25];
        eta_sum[7][26]  = eta_sum_out_tmp[7][26];
        eta_sum[7][27]  = eta_sum_out_tmp[7][27];
        eta_sum[7][28]  = eta_sum_out_tmp[7][28];
        eta_sum[7][29]  = eta_sum_out_tmp[7][29];
        eta_sum[7][30]  = eta_sum_out_tmp[7][30];
        eta_sum[7][31]  = eta_sum_out_tmp[7][31];
        eta_sum[7][32]  = eta_sum_out_tmp[7][32];
        eta_sum[7][33]  = eta_sum_out_tmp[7][33];
        eta_sum[7][34]  = eta_sum_out_tmp[7][34];
        eta_sum[7][35]  = eta_sum_out_tmp[7][35];
        eta_sum[7][36]  = eta_sum_out_tmp[7][36];
        eta_sum[7][37]  = eta_sum_out_tmp[7][37];
        eta_sum[7][38]  = eta_sum_out_tmp[7][38];
        eta_sum[7][39]  = eta_sum_out_tmp[7][39];
        eta_sum[7][40]  = eta_sum_out_tmp[7][40];
        eta_sum[7][41]  = eta_sum_out_tmp[7][41];
    end
 
endcase
end

if (chk_n_output_valid[0] & active_cols[8]) begin
case (curr_layer)
    0:begin 
        eta_sum[8][18]  = eta_sum_out_tmp[8][0];
        eta_sum[8][19]  = eta_sum_out_tmp[8][1];
        eta_sum[8][20]  = eta_sum_out_tmp[8][2];
        eta_sum[8][21]  = eta_sum_out_tmp[8][3];
        eta_sum[8][22]  = eta_sum_out_tmp[8][4];
        eta_sum[8][23]  = eta_sum_out_tmp[8][5];
        eta_sum[8][24]  = eta_sum_out_tmp[8][6];
        eta_sum[8][25]  = eta_sum_out_tmp[8][7];
        eta_sum[8][26]  = eta_sum_out_tmp[8][8];
        eta_sum[8][27]  = eta_sum_out_tmp[8][9];
        eta_sum[8][28]  = eta_sum_out_tmp[8][10];
        eta_sum[8][29]  = eta_sum_out_tmp[8][11];
        eta_sum[8][30]  = eta_sum_out_tmp[8][12];
        eta_sum[8][31]  = eta_sum_out_tmp[8][13];
        eta_sum[8][32]  = eta_sum_out_tmp[8][14];
        eta_sum[8][33]  = eta_sum_out_tmp[8][15];
        eta_sum[8][34]  = eta_sum_out_tmp[8][16];
        eta_sum[8][35]  = eta_sum_out_tmp[8][17];
        eta_sum[8][36]  = eta_sum_out_tmp[8][18];
        eta_sum[8][37]  = eta_sum_out_tmp[8][19];
        eta_sum[8][38]  = eta_sum_out_tmp[8][20];
        eta_sum[8][39]  = eta_sum_out_tmp[8][21];
        eta_sum[8][40]  = eta_sum_out_tmp[8][22];
        eta_sum[8][41]  = eta_sum_out_tmp[8][23];
        eta_sum[8][0]  = eta_sum_out_tmp[8][24];
        eta_sum[8][1]  = eta_sum_out_tmp[8][25];
        eta_sum[8][2]  = eta_sum_out_tmp[8][26];
        eta_sum[8][3]  = eta_sum_out_tmp[8][27];
        eta_sum[8][4]  = eta_sum_out_tmp[8][28];
        eta_sum[8][5]  = eta_sum_out_tmp[8][29];
        eta_sum[8][6]  = eta_sum_out_tmp[8][30];
        eta_sum[8][7]  = eta_sum_out_tmp[8][31];
        eta_sum[8][8]  = eta_sum_out_tmp[8][32];
        eta_sum[8][9]  = eta_sum_out_tmp[8][33];
        eta_sum[8][10]  = eta_sum_out_tmp[8][34];
        eta_sum[8][11]  = eta_sum_out_tmp[8][35];
        eta_sum[8][12]  = eta_sum_out_tmp[8][36];
        eta_sum[8][13]  = eta_sum_out_tmp[8][37];
        eta_sum[8][14]  = eta_sum_out_tmp[8][38];
        eta_sum[8][15]  = eta_sum_out_tmp[8][39];
        eta_sum[8][16]  = eta_sum_out_tmp[8][40];
        eta_sum[8][17]  = eta_sum_out_tmp[8][41];
    end
 
    1:begin 
        eta_sum[8][2]  = eta_sum_out_tmp[8][0];
        eta_sum[8][3]  = eta_sum_out_tmp[8][1];
        eta_sum[8][4]  = eta_sum_out_tmp[8][2];
        eta_sum[8][5]  = eta_sum_out_tmp[8][3];
        eta_sum[8][6]  = eta_sum_out_tmp[8][4];
        eta_sum[8][7]  = eta_sum_out_tmp[8][5];
        eta_sum[8][8]  = eta_sum_out_tmp[8][6];
        eta_sum[8][9]  = eta_sum_out_tmp[8][7];
        eta_sum[8][10]  = eta_sum_out_tmp[8][8];
        eta_sum[8][11]  = eta_sum_out_tmp[8][9];
        eta_sum[8][12]  = eta_sum_out_tmp[8][10];
        eta_sum[8][13]  = eta_sum_out_tmp[8][11];
        eta_sum[8][14]  = eta_sum_out_tmp[8][12];
        eta_sum[8][15]  = eta_sum_out_tmp[8][13];
        eta_sum[8][16]  = eta_sum_out_tmp[8][14];
        eta_sum[8][17]  = eta_sum_out_tmp[8][15];
        eta_sum[8][18]  = eta_sum_out_tmp[8][16];
        eta_sum[8][19]  = eta_sum_out_tmp[8][17];
        eta_sum[8][20]  = eta_sum_out_tmp[8][18];
        eta_sum[8][21]  = eta_sum_out_tmp[8][19];
        eta_sum[8][22]  = eta_sum_out_tmp[8][20];
        eta_sum[8][23]  = eta_sum_out_tmp[8][21];
        eta_sum[8][24]  = eta_sum_out_tmp[8][22];
        eta_sum[8][25]  = eta_sum_out_tmp[8][23];
        eta_sum[8][26]  = eta_sum_out_tmp[8][24];
        eta_sum[8][27]  = eta_sum_out_tmp[8][25];
        eta_sum[8][28]  = eta_sum_out_tmp[8][26];
        eta_sum[8][29]  = eta_sum_out_tmp[8][27];
        eta_sum[8][30]  = eta_sum_out_tmp[8][28];
        eta_sum[8][31]  = eta_sum_out_tmp[8][29];
        eta_sum[8][32]  = eta_sum_out_tmp[8][30];
        eta_sum[8][33]  = eta_sum_out_tmp[8][31];
        eta_sum[8][34]  = eta_sum_out_tmp[8][32];
        eta_sum[8][35]  = eta_sum_out_tmp[8][33];
        eta_sum[8][36]  = eta_sum_out_tmp[8][34];
        eta_sum[8][37]  = eta_sum_out_tmp[8][35];
        eta_sum[8][38]  = eta_sum_out_tmp[8][36];
        eta_sum[8][39]  = eta_sum_out_tmp[8][37];
        eta_sum[8][40]  = eta_sum_out_tmp[8][38];
        eta_sum[8][41]  = eta_sum_out_tmp[8][39];
        eta_sum[8][0]  = eta_sum_out_tmp[8][40];
        eta_sum[8][1]  = eta_sum_out_tmp[8][41];
    end
 
    2:begin 
        eta_sum[8][0]  = eta_sum_out_tmp[8][0];
        eta_sum[8][1]  = eta_sum_out_tmp[8][1];
        eta_sum[8][2]  = eta_sum_out_tmp[8][2];
        eta_sum[8][3]  = eta_sum_out_tmp[8][3];
        eta_sum[8][4]  = eta_sum_out_tmp[8][4];
        eta_sum[8][5]  = eta_sum_out_tmp[8][5];
        eta_sum[8][6]  = eta_sum_out_tmp[8][6];
        eta_sum[8][7]  = eta_sum_out_tmp[8][7];
        eta_sum[8][8]  = eta_sum_out_tmp[8][8];
        eta_sum[8][9]  = eta_sum_out_tmp[8][9];
        eta_sum[8][10]  = eta_sum_out_tmp[8][10];
        eta_sum[8][11]  = eta_sum_out_tmp[8][11];
        eta_sum[8][12]  = eta_sum_out_tmp[8][12];
        eta_sum[8][13]  = eta_sum_out_tmp[8][13];
        eta_sum[8][14]  = eta_sum_out_tmp[8][14];
        eta_sum[8][15]  = eta_sum_out_tmp[8][15];
        eta_sum[8][16]  = eta_sum_out_tmp[8][16];
        eta_sum[8][17]  = eta_sum_out_tmp[8][17];
        eta_sum[8][18]  = eta_sum_out_tmp[8][18];
        eta_sum[8][19]  = eta_sum_out_tmp[8][19];
        eta_sum[8][20]  = eta_sum_out_tmp[8][20];
        eta_sum[8][21]  = eta_sum_out_tmp[8][21];
        eta_sum[8][22]  = eta_sum_out_tmp[8][22];
        eta_sum[8][23]  = eta_sum_out_tmp[8][23];
        eta_sum[8][24]  = eta_sum_out_tmp[8][24];
        eta_sum[8][25]  = eta_sum_out_tmp[8][25];
        eta_sum[8][26]  = eta_sum_out_tmp[8][26];
        eta_sum[8][27]  = eta_sum_out_tmp[8][27];
        eta_sum[8][28]  = eta_sum_out_tmp[8][28];
        eta_sum[8][29]  = eta_sum_out_tmp[8][29];
        eta_sum[8][30]  = eta_sum_out_tmp[8][30];
        eta_sum[8][31]  = eta_sum_out_tmp[8][31];
        eta_sum[8][32]  = eta_sum_out_tmp[8][32];
        eta_sum[8][33]  = eta_sum_out_tmp[8][33];
        eta_sum[8][34]  = eta_sum_out_tmp[8][34];
        eta_sum[8][35]  = eta_sum_out_tmp[8][35];
        eta_sum[8][36]  = eta_sum_out_tmp[8][36];
        eta_sum[8][37]  = eta_sum_out_tmp[8][37];
        eta_sum[8][38]  = eta_sum_out_tmp[8][38];
        eta_sum[8][39]  = eta_sum_out_tmp[8][39];
        eta_sum[8][40]  = eta_sum_out_tmp[8][40];
        eta_sum[8][41]  = eta_sum_out_tmp[8][41];
    end
 
    3:begin 
        eta_sum[8][0]  = eta_sum_out_tmp[8][0];
        eta_sum[8][1]  = eta_sum_out_tmp[8][1];
        eta_sum[8][2]  = eta_sum_out_tmp[8][2];
        eta_sum[8][3]  = eta_sum_out_tmp[8][3];
        eta_sum[8][4]  = eta_sum_out_tmp[8][4];
        eta_sum[8][5]  = eta_sum_out_tmp[8][5];
        eta_sum[8][6]  = eta_sum_out_tmp[8][6];
        eta_sum[8][7]  = eta_sum_out_tmp[8][7];
        eta_sum[8][8]  = eta_sum_out_tmp[8][8];
        eta_sum[8][9]  = eta_sum_out_tmp[8][9];
        eta_sum[8][10]  = eta_sum_out_tmp[8][10];
        eta_sum[8][11]  = eta_sum_out_tmp[8][11];
        eta_sum[8][12]  = eta_sum_out_tmp[8][12];
        eta_sum[8][13]  = eta_sum_out_tmp[8][13];
        eta_sum[8][14]  = eta_sum_out_tmp[8][14];
        eta_sum[8][15]  = eta_sum_out_tmp[8][15];
        eta_sum[8][16]  = eta_sum_out_tmp[8][16];
        eta_sum[8][17]  = eta_sum_out_tmp[8][17];
        eta_sum[8][18]  = eta_sum_out_tmp[8][18];
        eta_sum[8][19]  = eta_sum_out_tmp[8][19];
        eta_sum[8][20]  = eta_sum_out_tmp[8][20];
        eta_sum[8][21]  = eta_sum_out_tmp[8][21];
        eta_sum[8][22]  = eta_sum_out_tmp[8][22];
        eta_sum[8][23]  = eta_sum_out_tmp[8][23];
        eta_sum[8][24]  = eta_sum_out_tmp[8][24];
        eta_sum[8][25]  = eta_sum_out_tmp[8][25];
        eta_sum[8][26]  = eta_sum_out_tmp[8][26];
        eta_sum[8][27]  = eta_sum_out_tmp[8][27];
        eta_sum[8][28]  = eta_sum_out_tmp[8][28];
        eta_sum[8][29]  = eta_sum_out_tmp[8][29];
        eta_sum[8][30]  = eta_sum_out_tmp[8][30];
        eta_sum[8][31]  = eta_sum_out_tmp[8][31];
        eta_sum[8][32]  = eta_sum_out_tmp[8][32];
        eta_sum[8][33]  = eta_sum_out_tmp[8][33];
        eta_sum[8][34]  = eta_sum_out_tmp[8][34];
        eta_sum[8][35]  = eta_sum_out_tmp[8][35];
        eta_sum[8][36]  = eta_sum_out_tmp[8][36];
        eta_sum[8][37]  = eta_sum_out_tmp[8][37];
        eta_sum[8][38]  = eta_sum_out_tmp[8][38];
        eta_sum[8][39]  = eta_sum_out_tmp[8][39];
        eta_sum[8][40]  = eta_sum_out_tmp[8][40];
        eta_sum[8][41]  = eta_sum_out_tmp[8][41];
    end
 
    4:begin 
        eta_sum[8][28]  = eta_sum_out_tmp[8][0];
        eta_sum[8][29]  = eta_sum_out_tmp[8][1];
        eta_sum[8][30]  = eta_sum_out_tmp[8][2];
        eta_sum[8][31]  = eta_sum_out_tmp[8][3];
        eta_sum[8][32]  = eta_sum_out_tmp[8][4];
        eta_sum[8][33]  = eta_sum_out_tmp[8][5];
        eta_sum[8][34]  = eta_sum_out_tmp[8][6];
        eta_sum[8][35]  = eta_sum_out_tmp[8][7];
        eta_sum[8][36]  = eta_sum_out_tmp[8][8];
        eta_sum[8][37]  = eta_sum_out_tmp[8][9];
        eta_sum[8][38]  = eta_sum_out_tmp[8][10];
        eta_sum[8][39]  = eta_sum_out_tmp[8][11];
        eta_sum[8][40]  = eta_sum_out_tmp[8][12];
        eta_sum[8][41]  = eta_sum_out_tmp[8][13];
        eta_sum[8][0]  = eta_sum_out_tmp[8][14];
        eta_sum[8][1]  = eta_sum_out_tmp[8][15];
        eta_sum[8][2]  = eta_sum_out_tmp[8][16];
        eta_sum[8][3]  = eta_sum_out_tmp[8][17];
        eta_sum[8][4]  = eta_sum_out_tmp[8][18];
        eta_sum[8][5]  = eta_sum_out_tmp[8][19];
        eta_sum[8][6]  = eta_sum_out_tmp[8][20];
        eta_sum[8][7]  = eta_sum_out_tmp[8][21];
        eta_sum[8][8]  = eta_sum_out_tmp[8][22];
        eta_sum[8][9]  = eta_sum_out_tmp[8][23];
        eta_sum[8][10]  = eta_sum_out_tmp[8][24];
        eta_sum[8][11]  = eta_sum_out_tmp[8][25];
        eta_sum[8][12]  = eta_sum_out_tmp[8][26];
        eta_sum[8][13]  = eta_sum_out_tmp[8][27];
        eta_sum[8][14]  = eta_sum_out_tmp[8][28];
        eta_sum[8][15]  = eta_sum_out_tmp[8][29];
        eta_sum[8][16]  = eta_sum_out_tmp[8][30];
        eta_sum[8][17]  = eta_sum_out_tmp[8][31];
        eta_sum[8][18]  = eta_sum_out_tmp[8][32];
        eta_sum[8][19]  = eta_sum_out_tmp[8][33];
        eta_sum[8][20]  = eta_sum_out_tmp[8][34];
        eta_sum[8][21]  = eta_sum_out_tmp[8][35];
        eta_sum[8][22]  = eta_sum_out_tmp[8][36];
        eta_sum[8][23]  = eta_sum_out_tmp[8][37];
        eta_sum[8][24]  = eta_sum_out_tmp[8][38];
        eta_sum[8][25]  = eta_sum_out_tmp[8][39];
        eta_sum[8][26]  = eta_sum_out_tmp[8][40];
        eta_sum[8][27]  = eta_sum_out_tmp[8][41];
    end
 
    5:begin 
        eta_sum[8][0]  = eta_sum_out_tmp[8][0];
        eta_sum[8][1]  = eta_sum_out_tmp[8][1];
        eta_sum[8][2]  = eta_sum_out_tmp[8][2];
        eta_sum[8][3]  = eta_sum_out_tmp[8][3];
        eta_sum[8][4]  = eta_sum_out_tmp[8][4];
        eta_sum[8][5]  = eta_sum_out_tmp[8][5];
        eta_sum[8][6]  = eta_sum_out_tmp[8][6];
        eta_sum[8][7]  = eta_sum_out_tmp[8][7];
        eta_sum[8][8]  = eta_sum_out_tmp[8][8];
        eta_sum[8][9]  = eta_sum_out_tmp[8][9];
        eta_sum[8][10]  = eta_sum_out_tmp[8][10];
        eta_sum[8][11]  = eta_sum_out_tmp[8][11];
        eta_sum[8][12]  = eta_sum_out_tmp[8][12];
        eta_sum[8][13]  = eta_sum_out_tmp[8][13];
        eta_sum[8][14]  = eta_sum_out_tmp[8][14];
        eta_sum[8][15]  = eta_sum_out_tmp[8][15];
        eta_sum[8][16]  = eta_sum_out_tmp[8][16];
        eta_sum[8][17]  = eta_sum_out_tmp[8][17];
        eta_sum[8][18]  = eta_sum_out_tmp[8][18];
        eta_sum[8][19]  = eta_sum_out_tmp[8][19];
        eta_sum[8][20]  = eta_sum_out_tmp[8][20];
        eta_sum[8][21]  = eta_sum_out_tmp[8][21];
        eta_sum[8][22]  = eta_sum_out_tmp[8][22];
        eta_sum[8][23]  = eta_sum_out_tmp[8][23];
        eta_sum[8][24]  = eta_sum_out_tmp[8][24];
        eta_sum[8][25]  = eta_sum_out_tmp[8][25];
        eta_sum[8][26]  = eta_sum_out_tmp[8][26];
        eta_sum[8][27]  = eta_sum_out_tmp[8][27];
        eta_sum[8][28]  = eta_sum_out_tmp[8][28];
        eta_sum[8][29]  = eta_sum_out_tmp[8][29];
        eta_sum[8][30]  = eta_sum_out_tmp[8][30];
        eta_sum[8][31]  = eta_sum_out_tmp[8][31];
        eta_sum[8][32]  = eta_sum_out_tmp[8][32];
        eta_sum[8][33]  = eta_sum_out_tmp[8][33];
        eta_sum[8][34]  = eta_sum_out_tmp[8][34];
        eta_sum[8][35]  = eta_sum_out_tmp[8][35];
        eta_sum[8][36]  = eta_sum_out_tmp[8][36];
        eta_sum[8][37]  = eta_sum_out_tmp[8][37];
        eta_sum[8][38]  = eta_sum_out_tmp[8][38];
        eta_sum[8][39]  = eta_sum_out_tmp[8][39];
        eta_sum[8][40]  = eta_sum_out_tmp[8][40];
        eta_sum[8][41]  = eta_sum_out_tmp[8][41];
    end
 
    6:begin 
        eta_sum[8][0]  = eta_sum_out_tmp[8][0];
        eta_sum[8][1]  = eta_sum_out_tmp[8][1];
        eta_sum[8][2]  = eta_sum_out_tmp[8][2];
        eta_sum[8][3]  = eta_sum_out_tmp[8][3];
        eta_sum[8][4]  = eta_sum_out_tmp[8][4];
        eta_sum[8][5]  = eta_sum_out_tmp[8][5];
        eta_sum[8][6]  = eta_sum_out_tmp[8][6];
        eta_sum[8][7]  = eta_sum_out_tmp[8][7];
        eta_sum[8][8]  = eta_sum_out_tmp[8][8];
        eta_sum[8][9]  = eta_sum_out_tmp[8][9];
        eta_sum[8][10]  = eta_sum_out_tmp[8][10];
        eta_sum[8][11]  = eta_sum_out_tmp[8][11];
        eta_sum[8][12]  = eta_sum_out_tmp[8][12];
        eta_sum[8][13]  = eta_sum_out_tmp[8][13];
        eta_sum[8][14]  = eta_sum_out_tmp[8][14];
        eta_sum[8][15]  = eta_sum_out_tmp[8][15];
        eta_sum[8][16]  = eta_sum_out_tmp[8][16];
        eta_sum[8][17]  = eta_sum_out_tmp[8][17];
        eta_sum[8][18]  = eta_sum_out_tmp[8][18];
        eta_sum[8][19]  = eta_sum_out_tmp[8][19];
        eta_sum[8][20]  = eta_sum_out_tmp[8][20];
        eta_sum[8][21]  = eta_sum_out_tmp[8][21];
        eta_sum[8][22]  = eta_sum_out_tmp[8][22];
        eta_sum[8][23]  = eta_sum_out_tmp[8][23];
        eta_sum[8][24]  = eta_sum_out_tmp[8][24];
        eta_sum[8][25]  = eta_sum_out_tmp[8][25];
        eta_sum[8][26]  = eta_sum_out_tmp[8][26];
        eta_sum[8][27]  = eta_sum_out_tmp[8][27];
        eta_sum[8][28]  = eta_sum_out_tmp[8][28];
        eta_sum[8][29]  = eta_sum_out_tmp[8][29];
        eta_sum[8][30]  = eta_sum_out_tmp[8][30];
        eta_sum[8][31]  = eta_sum_out_tmp[8][31];
        eta_sum[8][32]  = eta_sum_out_tmp[8][32];
        eta_sum[8][33]  = eta_sum_out_tmp[8][33];
        eta_sum[8][34]  = eta_sum_out_tmp[8][34];
        eta_sum[8][35]  = eta_sum_out_tmp[8][35];
        eta_sum[8][36]  = eta_sum_out_tmp[8][36];
        eta_sum[8][37]  = eta_sum_out_tmp[8][37];
        eta_sum[8][38]  = eta_sum_out_tmp[8][38];
        eta_sum[8][39]  = eta_sum_out_tmp[8][39];
        eta_sum[8][40]  = eta_sum_out_tmp[8][40];
        eta_sum[8][41]  = eta_sum_out_tmp[8][41];
    end
 
    7:begin 
        eta_sum[8][4]  = eta_sum_out_tmp[8][0];
        eta_sum[8][5]  = eta_sum_out_tmp[8][1];
        eta_sum[8][6]  = eta_sum_out_tmp[8][2];
        eta_sum[8][7]  = eta_sum_out_tmp[8][3];
        eta_sum[8][8]  = eta_sum_out_tmp[8][4];
        eta_sum[8][9]  = eta_sum_out_tmp[8][5];
        eta_sum[8][10]  = eta_sum_out_tmp[8][6];
        eta_sum[8][11]  = eta_sum_out_tmp[8][7];
        eta_sum[8][12]  = eta_sum_out_tmp[8][8];
        eta_sum[8][13]  = eta_sum_out_tmp[8][9];
        eta_sum[8][14]  = eta_sum_out_tmp[8][10];
        eta_sum[8][15]  = eta_sum_out_tmp[8][11];
        eta_sum[8][16]  = eta_sum_out_tmp[8][12];
        eta_sum[8][17]  = eta_sum_out_tmp[8][13];
        eta_sum[8][18]  = eta_sum_out_tmp[8][14];
        eta_sum[8][19]  = eta_sum_out_tmp[8][15];
        eta_sum[8][20]  = eta_sum_out_tmp[8][16];
        eta_sum[8][21]  = eta_sum_out_tmp[8][17];
        eta_sum[8][22]  = eta_sum_out_tmp[8][18];
        eta_sum[8][23]  = eta_sum_out_tmp[8][19];
        eta_sum[8][24]  = eta_sum_out_tmp[8][20];
        eta_sum[8][25]  = eta_sum_out_tmp[8][21];
        eta_sum[8][26]  = eta_sum_out_tmp[8][22];
        eta_sum[8][27]  = eta_sum_out_tmp[8][23];
        eta_sum[8][28]  = eta_sum_out_tmp[8][24];
        eta_sum[8][29]  = eta_sum_out_tmp[8][25];
        eta_sum[8][30]  = eta_sum_out_tmp[8][26];
        eta_sum[8][31]  = eta_sum_out_tmp[8][27];
        eta_sum[8][32]  = eta_sum_out_tmp[8][28];
        eta_sum[8][33]  = eta_sum_out_tmp[8][29];
        eta_sum[8][34]  = eta_sum_out_tmp[8][30];
        eta_sum[8][35]  = eta_sum_out_tmp[8][31];
        eta_sum[8][36]  = eta_sum_out_tmp[8][32];
        eta_sum[8][37]  = eta_sum_out_tmp[8][33];
        eta_sum[8][38]  = eta_sum_out_tmp[8][34];
        eta_sum[8][39]  = eta_sum_out_tmp[8][35];
        eta_sum[8][40]  = eta_sum_out_tmp[8][36];
        eta_sum[8][41]  = eta_sum_out_tmp[8][37];
        eta_sum[8][0]  = eta_sum_out_tmp[8][38];
        eta_sum[8][1]  = eta_sum_out_tmp[8][39];
        eta_sum[8][2]  = eta_sum_out_tmp[8][40];
        eta_sum[8][3]  = eta_sum_out_tmp[8][41];
    end
 
endcase
end

if (chk_n_output_valid[0] & active_cols[9]) begin
case (curr_layer)
    0:begin 
        eta_sum[9][0]  = eta_sum_out_tmp[9][0];
        eta_sum[9][1]  = eta_sum_out_tmp[9][1];
        eta_sum[9][2]  = eta_sum_out_tmp[9][2];
        eta_sum[9][3]  = eta_sum_out_tmp[9][3];
        eta_sum[9][4]  = eta_sum_out_tmp[9][4];
        eta_sum[9][5]  = eta_sum_out_tmp[9][5];
        eta_sum[9][6]  = eta_sum_out_tmp[9][6];
        eta_sum[9][7]  = eta_sum_out_tmp[9][7];
        eta_sum[9][8]  = eta_sum_out_tmp[9][8];
        eta_sum[9][9]  = eta_sum_out_tmp[9][9];
        eta_sum[9][10]  = eta_sum_out_tmp[9][10];
        eta_sum[9][11]  = eta_sum_out_tmp[9][11];
        eta_sum[9][12]  = eta_sum_out_tmp[9][12];
        eta_sum[9][13]  = eta_sum_out_tmp[9][13];
        eta_sum[9][14]  = eta_sum_out_tmp[9][14];
        eta_sum[9][15]  = eta_sum_out_tmp[9][15];
        eta_sum[9][16]  = eta_sum_out_tmp[9][16];
        eta_sum[9][17]  = eta_sum_out_tmp[9][17];
        eta_sum[9][18]  = eta_sum_out_tmp[9][18];
        eta_sum[9][19]  = eta_sum_out_tmp[9][19];
        eta_sum[9][20]  = eta_sum_out_tmp[9][20];
        eta_sum[9][21]  = eta_sum_out_tmp[9][21];
        eta_sum[9][22]  = eta_sum_out_tmp[9][22];
        eta_sum[9][23]  = eta_sum_out_tmp[9][23];
        eta_sum[9][24]  = eta_sum_out_tmp[9][24];
        eta_sum[9][25]  = eta_sum_out_tmp[9][25];
        eta_sum[9][26]  = eta_sum_out_tmp[9][26];
        eta_sum[9][27]  = eta_sum_out_tmp[9][27];
        eta_sum[9][28]  = eta_sum_out_tmp[9][28];
        eta_sum[9][29]  = eta_sum_out_tmp[9][29];
        eta_sum[9][30]  = eta_sum_out_tmp[9][30];
        eta_sum[9][31]  = eta_sum_out_tmp[9][31];
        eta_sum[9][32]  = eta_sum_out_tmp[9][32];
        eta_sum[9][33]  = eta_sum_out_tmp[9][33];
        eta_sum[9][34]  = eta_sum_out_tmp[9][34];
        eta_sum[9][35]  = eta_sum_out_tmp[9][35];
        eta_sum[9][36]  = eta_sum_out_tmp[9][36];
        eta_sum[9][37]  = eta_sum_out_tmp[9][37];
        eta_sum[9][38]  = eta_sum_out_tmp[9][38];
        eta_sum[9][39]  = eta_sum_out_tmp[9][39];
        eta_sum[9][40]  = eta_sum_out_tmp[9][40];
        eta_sum[9][41]  = eta_sum_out_tmp[9][41];
    end
 
    1:begin 
        eta_sum[9][1]  = eta_sum_out_tmp[9][0];
        eta_sum[9][2]  = eta_sum_out_tmp[9][1];
        eta_sum[9][3]  = eta_sum_out_tmp[9][2];
        eta_sum[9][4]  = eta_sum_out_tmp[9][3];
        eta_sum[9][5]  = eta_sum_out_tmp[9][4];
        eta_sum[9][6]  = eta_sum_out_tmp[9][5];
        eta_sum[9][7]  = eta_sum_out_tmp[9][6];
        eta_sum[9][8]  = eta_sum_out_tmp[9][7];
        eta_sum[9][9]  = eta_sum_out_tmp[9][8];
        eta_sum[9][10]  = eta_sum_out_tmp[9][9];
        eta_sum[9][11]  = eta_sum_out_tmp[9][10];
        eta_sum[9][12]  = eta_sum_out_tmp[9][11];
        eta_sum[9][13]  = eta_sum_out_tmp[9][12];
        eta_sum[9][14]  = eta_sum_out_tmp[9][13];
        eta_sum[9][15]  = eta_sum_out_tmp[9][14];
        eta_sum[9][16]  = eta_sum_out_tmp[9][15];
        eta_sum[9][17]  = eta_sum_out_tmp[9][16];
        eta_sum[9][18]  = eta_sum_out_tmp[9][17];
        eta_sum[9][19]  = eta_sum_out_tmp[9][18];
        eta_sum[9][20]  = eta_sum_out_tmp[9][19];
        eta_sum[9][21]  = eta_sum_out_tmp[9][20];
        eta_sum[9][22]  = eta_sum_out_tmp[9][21];
        eta_sum[9][23]  = eta_sum_out_tmp[9][22];
        eta_sum[9][24]  = eta_sum_out_tmp[9][23];
        eta_sum[9][25]  = eta_sum_out_tmp[9][24];
        eta_sum[9][26]  = eta_sum_out_tmp[9][25];
        eta_sum[9][27]  = eta_sum_out_tmp[9][26];
        eta_sum[9][28]  = eta_sum_out_tmp[9][27];
        eta_sum[9][29]  = eta_sum_out_tmp[9][28];
        eta_sum[9][30]  = eta_sum_out_tmp[9][29];
        eta_sum[9][31]  = eta_sum_out_tmp[9][30];
        eta_sum[9][32]  = eta_sum_out_tmp[9][31];
        eta_sum[9][33]  = eta_sum_out_tmp[9][32];
        eta_sum[9][34]  = eta_sum_out_tmp[9][33];
        eta_sum[9][35]  = eta_sum_out_tmp[9][34];
        eta_sum[9][36]  = eta_sum_out_tmp[9][35];
        eta_sum[9][37]  = eta_sum_out_tmp[9][36];
        eta_sum[9][38]  = eta_sum_out_tmp[9][37];
        eta_sum[9][39]  = eta_sum_out_tmp[9][38];
        eta_sum[9][40]  = eta_sum_out_tmp[9][39];
        eta_sum[9][41]  = eta_sum_out_tmp[9][40];
        eta_sum[9][0]  = eta_sum_out_tmp[9][41];
    end
 
    2:begin 
        eta_sum[9][10]  = eta_sum_out_tmp[9][0];
        eta_sum[9][11]  = eta_sum_out_tmp[9][1];
        eta_sum[9][12]  = eta_sum_out_tmp[9][2];
        eta_sum[9][13]  = eta_sum_out_tmp[9][3];
        eta_sum[9][14]  = eta_sum_out_tmp[9][4];
        eta_sum[9][15]  = eta_sum_out_tmp[9][5];
        eta_sum[9][16]  = eta_sum_out_tmp[9][6];
        eta_sum[9][17]  = eta_sum_out_tmp[9][7];
        eta_sum[9][18]  = eta_sum_out_tmp[9][8];
        eta_sum[9][19]  = eta_sum_out_tmp[9][9];
        eta_sum[9][20]  = eta_sum_out_tmp[9][10];
        eta_sum[9][21]  = eta_sum_out_tmp[9][11];
        eta_sum[9][22]  = eta_sum_out_tmp[9][12];
        eta_sum[9][23]  = eta_sum_out_tmp[9][13];
        eta_sum[9][24]  = eta_sum_out_tmp[9][14];
        eta_sum[9][25]  = eta_sum_out_tmp[9][15];
        eta_sum[9][26]  = eta_sum_out_tmp[9][16];
        eta_sum[9][27]  = eta_sum_out_tmp[9][17];
        eta_sum[9][28]  = eta_sum_out_tmp[9][18];
        eta_sum[9][29]  = eta_sum_out_tmp[9][19];
        eta_sum[9][30]  = eta_sum_out_tmp[9][20];
        eta_sum[9][31]  = eta_sum_out_tmp[9][21];
        eta_sum[9][32]  = eta_sum_out_tmp[9][22];
        eta_sum[9][33]  = eta_sum_out_tmp[9][23];
        eta_sum[9][34]  = eta_sum_out_tmp[9][24];
        eta_sum[9][35]  = eta_sum_out_tmp[9][25];
        eta_sum[9][36]  = eta_sum_out_tmp[9][26];
        eta_sum[9][37]  = eta_sum_out_tmp[9][27];
        eta_sum[9][38]  = eta_sum_out_tmp[9][28];
        eta_sum[9][39]  = eta_sum_out_tmp[9][29];
        eta_sum[9][40]  = eta_sum_out_tmp[9][30];
        eta_sum[9][41]  = eta_sum_out_tmp[9][31];
        eta_sum[9][0]  = eta_sum_out_tmp[9][32];
        eta_sum[9][1]  = eta_sum_out_tmp[9][33];
        eta_sum[9][2]  = eta_sum_out_tmp[9][34];
        eta_sum[9][3]  = eta_sum_out_tmp[9][35];
        eta_sum[9][4]  = eta_sum_out_tmp[9][36];
        eta_sum[9][5]  = eta_sum_out_tmp[9][37];
        eta_sum[9][6]  = eta_sum_out_tmp[9][38];
        eta_sum[9][7]  = eta_sum_out_tmp[9][39];
        eta_sum[9][8]  = eta_sum_out_tmp[9][40];
        eta_sum[9][9]  = eta_sum_out_tmp[9][41];
    end
 
    3:begin 
        eta_sum[9][0]  = eta_sum_out_tmp[9][0];
        eta_sum[9][1]  = eta_sum_out_tmp[9][1];
        eta_sum[9][2]  = eta_sum_out_tmp[9][2];
        eta_sum[9][3]  = eta_sum_out_tmp[9][3];
        eta_sum[9][4]  = eta_sum_out_tmp[9][4];
        eta_sum[9][5]  = eta_sum_out_tmp[9][5];
        eta_sum[9][6]  = eta_sum_out_tmp[9][6];
        eta_sum[9][7]  = eta_sum_out_tmp[9][7];
        eta_sum[9][8]  = eta_sum_out_tmp[9][8];
        eta_sum[9][9]  = eta_sum_out_tmp[9][9];
        eta_sum[9][10]  = eta_sum_out_tmp[9][10];
        eta_sum[9][11]  = eta_sum_out_tmp[9][11];
        eta_sum[9][12]  = eta_sum_out_tmp[9][12];
        eta_sum[9][13]  = eta_sum_out_tmp[9][13];
        eta_sum[9][14]  = eta_sum_out_tmp[9][14];
        eta_sum[9][15]  = eta_sum_out_tmp[9][15];
        eta_sum[9][16]  = eta_sum_out_tmp[9][16];
        eta_sum[9][17]  = eta_sum_out_tmp[9][17];
        eta_sum[9][18]  = eta_sum_out_tmp[9][18];
        eta_sum[9][19]  = eta_sum_out_tmp[9][19];
        eta_sum[9][20]  = eta_sum_out_tmp[9][20];
        eta_sum[9][21]  = eta_sum_out_tmp[9][21];
        eta_sum[9][22]  = eta_sum_out_tmp[9][22];
        eta_sum[9][23]  = eta_sum_out_tmp[9][23];
        eta_sum[9][24]  = eta_sum_out_tmp[9][24];
        eta_sum[9][25]  = eta_sum_out_tmp[9][25];
        eta_sum[9][26]  = eta_sum_out_tmp[9][26];
        eta_sum[9][27]  = eta_sum_out_tmp[9][27];
        eta_sum[9][28]  = eta_sum_out_tmp[9][28];
        eta_sum[9][29]  = eta_sum_out_tmp[9][29];
        eta_sum[9][30]  = eta_sum_out_tmp[9][30];
        eta_sum[9][31]  = eta_sum_out_tmp[9][31];
        eta_sum[9][32]  = eta_sum_out_tmp[9][32];
        eta_sum[9][33]  = eta_sum_out_tmp[9][33];
        eta_sum[9][34]  = eta_sum_out_tmp[9][34];
        eta_sum[9][35]  = eta_sum_out_tmp[9][35];
        eta_sum[9][36]  = eta_sum_out_tmp[9][36];
        eta_sum[9][37]  = eta_sum_out_tmp[9][37];
        eta_sum[9][38]  = eta_sum_out_tmp[9][38];
        eta_sum[9][39]  = eta_sum_out_tmp[9][39];
        eta_sum[9][40]  = eta_sum_out_tmp[9][40];
        eta_sum[9][41]  = eta_sum_out_tmp[9][41];
    end
 
    4:begin 
        eta_sum[9][0]  = eta_sum_out_tmp[9][0];
        eta_sum[9][1]  = eta_sum_out_tmp[9][1];
        eta_sum[9][2]  = eta_sum_out_tmp[9][2];
        eta_sum[9][3]  = eta_sum_out_tmp[9][3];
        eta_sum[9][4]  = eta_sum_out_tmp[9][4];
        eta_sum[9][5]  = eta_sum_out_tmp[9][5];
        eta_sum[9][6]  = eta_sum_out_tmp[9][6];
        eta_sum[9][7]  = eta_sum_out_tmp[9][7];
        eta_sum[9][8]  = eta_sum_out_tmp[9][8];
        eta_sum[9][9]  = eta_sum_out_tmp[9][9];
        eta_sum[9][10]  = eta_sum_out_tmp[9][10];
        eta_sum[9][11]  = eta_sum_out_tmp[9][11];
        eta_sum[9][12]  = eta_sum_out_tmp[9][12];
        eta_sum[9][13]  = eta_sum_out_tmp[9][13];
        eta_sum[9][14]  = eta_sum_out_tmp[9][14];
        eta_sum[9][15]  = eta_sum_out_tmp[9][15];
        eta_sum[9][16]  = eta_sum_out_tmp[9][16];
        eta_sum[9][17]  = eta_sum_out_tmp[9][17];
        eta_sum[9][18]  = eta_sum_out_tmp[9][18];
        eta_sum[9][19]  = eta_sum_out_tmp[9][19];
        eta_sum[9][20]  = eta_sum_out_tmp[9][20];
        eta_sum[9][21]  = eta_sum_out_tmp[9][21];
        eta_sum[9][22]  = eta_sum_out_tmp[9][22];
        eta_sum[9][23]  = eta_sum_out_tmp[9][23];
        eta_sum[9][24]  = eta_sum_out_tmp[9][24];
        eta_sum[9][25]  = eta_sum_out_tmp[9][25];
        eta_sum[9][26]  = eta_sum_out_tmp[9][26];
        eta_sum[9][27]  = eta_sum_out_tmp[9][27];
        eta_sum[9][28]  = eta_sum_out_tmp[9][28];
        eta_sum[9][29]  = eta_sum_out_tmp[9][29];
        eta_sum[9][30]  = eta_sum_out_tmp[9][30];
        eta_sum[9][31]  = eta_sum_out_tmp[9][31];
        eta_sum[9][32]  = eta_sum_out_tmp[9][32];
        eta_sum[9][33]  = eta_sum_out_tmp[9][33];
        eta_sum[9][34]  = eta_sum_out_tmp[9][34];
        eta_sum[9][35]  = eta_sum_out_tmp[9][35];
        eta_sum[9][36]  = eta_sum_out_tmp[9][36];
        eta_sum[9][37]  = eta_sum_out_tmp[9][37];
        eta_sum[9][38]  = eta_sum_out_tmp[9][38];
        eta_sum[9][39]  = eta_sum_out_tmp[9][39];
        eta_sum[9][40]  = eta_sum_out_tmp[9][40];
        eta_sum[9][41]  = eta_sum_out_tmp[9][41];
    end
 
    5:begin 
        eta_sum[9][28]  = eta_sum_out_tmp[9][0];
        eta_sum[9][29]  = eta_sum_out_tmp[9][1];
        eta_sum[9][30]  = eta_sum_out_tmp[9][2];
        eta_sum[9][31]  = eta_sum_out_tmp[9][3];
        eta_sum[9][32]  = eta_sum_out_tmp[9][4];
        eta_sum[9][33]  = eta_sum_out_tmp[9][5];
        eta_sum[9][34]  = eta_sum_out_tmp[9][6];
        eta_sum[9][35]  = eta_sum_out_tmp[9][7];
        eta_sum[9][36]  = eta_sum_out_tmp[9][8];
        eta_sum[9][37]  = eta_sum_out_tmp[9][9];
        eta_sum[9][38]  = eta_sum_out_tmp[9][10];
        eta_sum[9][39]  = eta_sum_out_tmp[9][11];
        eta_sum[9][40]  = eta_sum_out_tmp[9][12];
        eta_sum[9][41]  = eta_sum_out_tmp[9][13];
        eta_sum[9][0]  = eta_sum_out_tmp[9][14];
        eta_sum[9][1]  = eta_sum_out_tmp[9][15];
        eta_sum[9][2]  = eta_sum_out_tmp[9][16];
        eta_sum[9][3]  = eta_sum_out_tmp[9][17];
        eta_sum[9][4]  = eta_sum_out_tmp[9][18];
        eta_sum[9][5]  = eta_sum_out_tmp[9][19];
        eta_sum[9][6]  = eta_sum_out_tmp[9][20];
        eta_sum[9][7]  = eta_sum_out_tmp[9][21];
        eta_sum[9][8]  = eta_sum_out_tmp[9][22];
        eta_sum[9][9]  = eta_sum_out_tmp[9][23];
        eta_sum[9][10]  = eta_sum_out_tmp[9][24];
        eta_sum[9][11]  = eta_sum_out_tmp[9][25];
        eta_sum[9][12]  = eta_sum_out_tmp[9][26];
        eta_sum[9][13]  = eta_sum_out_tmp[9][27];
        eta_sum[9][14]  = eta_sum_out_tmp[9][28];
        eta_sum[9][15]  = eta_sum_out_tmp[9][29];
        eta_sum[9][16]  = eta_sum_out_tmp[9][30];
        eta_sum[9][17]  = eta_sum_out_tmp[9][31];
        eta_sum[9][18]  = eta_sum_out_tmp[9][32];
        eta_sum[9][19]  = eta_sum_out_tmp[9][33];
        eta_sum[9][20]  = eta_sum_out_tmp[9][34];
        eta_sum[9][21]  = eta_sum_out_tmp[9][35];
        eta_sum[9][22]  = eta_sum_out_tmp[9][36];
        eta_sum[9][23]  = eta_sum_out_tmp[9][37];
        eta_sum[9][24]  = eta_sum_out_tmp[9][38];
        eta_sum[9][25]  = eta_sum_out_tmp[9][39];
        eta_sum[9][26]  = eta_sum_out_tmp[9][40];
        eta_sum[9][27]  = eta_sum_out_tmp[9][41];
    end
 
    6:begin 
        eta_sum[9][0]  = eta_sum_out_tmp[9][0];
        eta_sum[9][1]  = eta_sum_out_tmp[9][1];
        eta_sum[9][2]  = eta_sum_out_tmp[9][2];
        eta_sum[9][3]  = eta_sum_out_tmp[9][3];
        eta_sum[9][4]  = eta_sum_out_tmp[9][4];
        eta_sum[9][5]  = eta_sum_out_tmp[9][5];
        eta_sum[9][6]  = eta_sum_out_tmp[9][6];
        eta_sum[9][7]  = eta_sum_out_tmp[9][7];
        eta_sum[9][8]  = eta_sum_out_tmp[9][8];
        eta_sum[9][9]  = eta_sum_out_tmp[9][9];
        eta_sum[9][10]  = eta_sum_out_tmp[9][10];
        eta_sum[9][11]  = eta_sum_out_tmp[9][11];
        eta_sum[9][12]  = eta_sum_out_tmp[9][12];
        eta_sum[9][13]  = eta_sum_out_tmp[9][13];
        eta_sum[9][14]  = eta_sum_out_tmp[9][14];
        eta_sum[9][15]  = eta_sum_out_tmp[9][15];
        eta_sum[9][16]  = eta_sum_out_tmp[9][16];
        eta_sum[9][17]  = eta_sum_out_tmp[9][17];
        eta_sum[9][18]  = eta_sum_out_tmp[9][18];
        eta_sum[9][19]  = eta_sum_out_tmp[9][19];
        eta_sum[9][20]  = eta_sum_out_tmp[9][20];
        eta_sum[9][21]  = eta_sum_out_tmp[9][21];
        eta_sum[9][22]  = eta_sum_out_tmp[9][22];
        eta_sum[9][23]  = eta_sum_out_tmp[9][23];
        eta_sum[9][24]  = eta_sum_out_tmp[9][24];
        eta_sum[9][25]  = eta_sum_out_tmp[9][25];
        eta_sum[9][26]  = eta_sum_out_tmp[9][26];
        eta_sum[9][27]  = eta_sum_out_tmp[9][27];
        eta_sum[9][28]  = eta_sum_out_tmp[9][28];
        eta_sum[9][29]  = eta_sum_out_tmp[9][29];
        eta_sum[9][30]  = eta_sum_out_tmp[9][30];
        eta_sum[9][31]  = eta_sum_out_tmp[9][31];
        eta_sum[9][32]  = eta_sum_out_tmp[9][32];
        eta_sum[9][33]  = eta_sum_out_tmp[9][33];
        eta_sum[9][34]  = eta_sum_out_tmp[9][34];
        eta_sum[9][35]  = eta_sum_out_tmp[9][35];
        eta_sum[9][36]  = eta_sum_out_tmp[9][36];
        eta_sum[9][37]  = eta_sum_out_tmp[9][37];
        eta_sum[9][38]  = eta_sum_out_tmp[9][38];
        eta_sum[9][39]  = eta_sum_out_tmp[9][39];
        eta_sum[9][40]  = eta_sum_out_tmp[9][40];
        eta_sum[9][41]  = eta_sum_out_tmp[9][41];
    end
 
    7:begin 
        eta_sum[9][0]  = eta_sum_out_tmp[9][0];
        eta_sum[9][1]  = eta_sum_out_tmp[9][1];
        eta_sum[9][2]  = eta_sum_out_tmp[9][2];
        eta_sum[9][3]  = eta_sum_out_tmp[9][3];
        eta_sum[9][4]  = eta_sum_out_tmp[9][4];
        eta_sum[9][5]  = eta_sum_out_tmp[9][5];
        eta_sum[9][6]  = eta_sum_out_tmp[9][6];
        eta_sum[9][7]  = eta_sum_out_tmp[9][7];
        eta_sum[9][8]  = eta_sum_out_tmp[9][8];
        eta_sum[9][9]  = eta_sum_out_tmp[9][9];
        eta_sum[9][10]  = eta_sum_out_tmp[9][10];
        eta_sum[9][11]  = eta_sum_out_tmp[9][11];
        eta_sum[9][12]  = eta_sum_out_tmp[9][12];
        eta_sum[9][13]  = eta_sum_out_tmp[9][13];
        eta_sum[9][14]  = eta_sum_out_tmp[9][14];
        eta_sum[9][15]  = eta_sum_out_tmp[9][15];
        eta_sum[9][16]  = eta_sum_out_tmp[9][16];
        eta_sum[9][17]  = eta_sum_out_tmp[9][17];
        eta_sum[9][18]  = eta_sum_out_tmp[9][18];
        eta_sum[9][19]  = eta_sum_out_tmp[9][19];
        eta_sum[9][20]  = eta_sum_out_tmp[9][20];
        eta_sum[9][21]  = eta_sum_out_tmp[9][21];
        eta_sum[9][22]  = eta_sum_out_tmp[9][22];
        eta_sum[9][23]  = eta_sum_out_tmp[9][23];
        eta_sum[9][24]  = eta_sum_out_tmp[9][24];
        eta_sum[9][25]  = eta_sum_out_tmp[9][25];
        eta_sum[9][26]  = eta_sum_out_tmp[9][26];
        eta_sum[9][27]  = eta_sum_out_tmp[9][27];
        eta_sum[9][28]  = eta_sum_out_tmp[9][28];
        eta_sum[9][29]  = eta_sum_out_tmp[9][29];
        eta_sum[9][30]  = eta_sum_out_tmp[9][30];
        eta_sum[9][31]  = eta_sum_out_tmp[9][31];
        eta_sum[9][32]  = eta_sum_out_tmp[9][32];
        eta_sum[9][33]  = eta_sum_out_tmp[9][33];
        eta_sum[9][34]  = eta_sum_out_tmp[9][34];
        eta_sum[9][35]  = eta_sum_out_tmp[9][35];
        eta_sum[9][36]  = eta_sum_out_tmp[9][36];
        eta_sum[9][37]  = eta_sum_out_tmp[9][37];
        eta_sum[9][38]  = eta_sum_out_tmp[9][38];
        eta_sum[9][39]  = eta_sum_out_tmp[9][39];
        eta_sum[9][40]  = eta_sum_out_tmp[9][40];
        eta_sum[9][41]  = eta_sum_out_tmp[9][41];
    end
 
endcase
end

if (chk_n_output_valid[0] & active_cols[10]) begin
case (curr_layer)
    0:begin 
        eta_sum[10][0]  = eta_sum_out_tmp[10][0];
        eta_sum[10][1]  = eta_sum_out_tmp[10][1];
        eta_sum[10][2]  = eta_sum_out_tmp[10][2];
        eta_sum[10][3]  = eta_sum_out_tmp[10][3];
        eta_sum[10][4]  = eta_sum_out_tmp[10][4];
        eta_sum[10][5]  = eta_sum_out_tmp[10][5];
        eta_sum[10][6]  = eta_sum_out_tmp[10][6];
        eta_sum[10][7]  = eta_sum_out_tmp[10][7];
        eta_sum[10][8]  = eta_sum_out_tmp[10][8];
        eta_sum[10][9]  = eta_sum_out_tmp[10][9];
        eta_sum[10][10]  = eta_sum_out_tmp[10][10];
        eta_sum[10][11]  = eta_sum_out_tmp[10][11];
        eta_sum[10][12]  = eta_sum_out_tmp[10][12];
        eta_sum[10][13]  = eta_sum_out_tmp[10][13];
        eta_sum[10][14]  = eta_sum_out_tmp[10][14];
        eta_sum[10][15]  = eta_sum_out_tmp[10][15];
        eta_sum[10][16]  = eta_sum_out_tmp[10][16];
        eta_sum[10][17]  = eta_sum_out_tmp[10][17];
        eta_sum[10][18]  = eta_sum_out_tmp[10][18];
        eta_sum[10][19]  = eta_sum_out_tmp[10][19];
        eta_sum[10][20]  = eta_sum_out_tmp[10][20];
        eta_sum[10][21]  = eta_sum_out_tmp[10][21];
        eta_sum[10][22]  = eta_sum_out_tmp[10][22];
        eta_sum[10][23]  = eta_sum_out_tmp[10][23];
        eta_sum[10][24]  = eta_sum_out_tmp[10][24];
        eta_sum[10][25]  = eta_sum_out_tmp[10][25];
        eta_sum[10][26]  = eta_sum_out_tmp[10][26];
        eta_sum[10][27]  = eta_sum_out_tmp[10][27];
        eta_sum[10][28]  = eta_sum_out_tmp[10][28];
        eta_sum[10][29]  = eta_sum_out_tmp[10][29];
        eta_sum[10][30]  = eta_sum_out_tmp[10][30];
        eta_sum[10][31]  = eta_sum_out_tmp[10][31];
        eta_sum[10][32]  = eta_sum_out_tmp[10][32];
        eta_sum[10][33]  = eta_sum_out_tmp[10][33];
        eta_sum[10][34]  = eta_sum_out_tmp[10][34];
        eta_sum[10][35]  = eta_sum_out_tmp[10][35];
        eta_sum[10][36]  = eta_sum_out_tmp[10][36];
        eta_sum[10][37]  = eta_sum_out_tmp[10][37];
        eta_sum[10][38]  = eta_sum_out_tmp[10][38];
        eta_sum[10][39]  = eta_sum_out_tmp[10][39];
        eta_sum[10][40]  = eta_sum_out_tmp[10][40];
        eta_sum[10][41]  = eta_sum_out_tmp[10][41];
    end
 
    1:begin 
        eta_sum[10][0]  = eta_sum_out_tmp[10][0];
        eta_sum[10][1]  = eta_sum_out_tmp[10][1];
        eta_sum[10][2]  = eta_sum_out_tmp[10][2];
        eta_sum[10][3]  = eta_sum_out_tmp[10][3];
        eta_sum[10][4]  = eta_sum_out_tmp[10][4];
        eta_sum[10][5]  = eta_sum_out_tmp[10][5];
        eta_sum[10][6]  = eta_sum_out_tmp[10][6];
        eta_sum[10][7]  = eta_sum_out_tmp[10][7];
        eta_sum[10][8]  = eta_sum_out_tmp[10][8];
        eta_sum[10][9]  = eta_sum_out_tmp[10][9];
        eta_sum[10][10]  = eta_sum_out_tmp[10][10];
        eta_sum[10][11]  = eta_sum_out_tmp[10][11];
        eta_sum[10][12]  = eta_sum_out_tmp[10][12];
        eta_sum[10][13]  = eta_sum_out_tmp[10][13];
        eta_sum[10][14]  = eta_sum_out_tmp[10][14];
        eta_sum[10][15]  = eta_sum_out_tmp[10][15];
        eta_sum[10][16]  = eta_sum_out_tmp[10][16];
        eta_sum[10][17]  = eta_sum_out_tmp[10][17];
        eta_sum[10][18]  = eta_sum_out_tmp[10][18];
        eta_sum[10][19]  = eta_sum_out_tmp[10][19];
        eta_sum[10][20]  = eta_sum_out_tmp[10][20];
        eta_sum[10][21]  = eta_sum_out_tmp[10][21];
        eta_sum[10][22]  = eta_sum_out_tmp[10][22];
        eta_sum[10][23]  = eta_sum_out_tmp[10][23];
        eta_sum[10][24]  = eta_sum_out_tmp[10][24];
        eta_sum[10][25]  = eta_sum_out_tmp[10][25];
        eta_sum[10][26]  = eta_sum_out_tmp[10][26];
        eta_sum[10][27]  = eta_sum_out_tmp[10][27];
        eta_sum[10][28]  = eta_sum_out_tmp[10][28];
        eta_sum[10][29]  = eta_sum_out_tmp[10][29];
        eta_sum[10][30]  = eta_sum_out_tmp[10][30];
        eta_sum[10][31]  = eta_sum_out_tmp[10][31];
        eta_sum[10][32]  = eta_sum_out_tmp[10][32];
        eta_sum[10][33]  = eta_sum_out_tmp[10][33];
        eta_sum[10][34]  = eta_sum_out_tmp[10][34];
        eta_sum[10][35]  = eta_sum_out_tmp[10][35];
        eta_sum[10][36]  = eta_sum_out_tmp[10][36];
        eta_sum[10][37]  = eta_sum_out_tmp[10][37];
        eta_sum[10][38]  = eta_sum_out_tmp[10][38];
        eta_sum[10][39]  = eta_sum_out_tmp[10][39];
        eta_sum[10][40]  = eta_sum_out_tmp[10][40];
        eta_sum[10][41]  = eta_sum_out_tmp[10][41];
    end
 
    2:begin 
        eta_sum[10][41]  = eta_sum_out_tmp[10][0];
        eta_sum[10][0]  = eta_sum_out_tmp[10][1];
        eta_sum[10][1]  = eta_sum_out_tmp[10][2];
        eta_sum[10][2]  = eta_sum_out_tmp[10][3];
        eta_sum[10][3]  = eta_sum_out_tmp[10][4];
        eta_sum[10][4]  = eta_sum_out_tmp[10][5];
        eta_sum[10][5]  = eta_sum_out_tmp[10][6];
        eta_sum[10][6]  = eta_sum_out_tmp[10][7];
        eta_sum[10][7]  = eta_sum_out_tmp[10][8];
        eta_sum[10][8]  = eta_sum_out_tmp[10][9];
        eta_sum[10][9]  = eta_sum_out_tmp[10][10];
        eta_sum[10][10]  = eta_sum_out_tmp[10][11];
        eta_sum[10][11]  = eta_sum_out_tmp[10][12];
        eta_sum[10][12]  = eta_sum_out_tmp[10][13];
        eta_sum[10][13]  = eta_sum_out_tmp[10][14];
        eta_sum[10][14]  = eta_sum_out_tmp[10][15];
        eta_sum[10][15]  = eta_sum_out_tmp[10][16];
        eta_sum[10][16]  = eta_sum_out_tmp[10][17];
        eta_sum[10][17]  = eta_sum_out_tmp[10][18];
        eta_sum[10][18]  = eta_sum_out_tmp[10][19];
        eta_sum[10][19]  = eta_sum_out_tmp[10][20];
        eta_sum[10][20]  = eta_sum_out_tmp[10][21];
        eta_sum[10][21]  = eta_sum_out_tmp[10][22];
        eta_sum[10][22]  = eta_sum_out_tmp[10][23];
        eta_sum[10][23]  = eta_sum_out_tmp[10][24];
        eta_sum[10][24]  = eta_sum_out_tmp[10][25];
        eta_sum[10][25]  = eta_sum_out_tmp[10][26];
        eta_sum[10][26]  = eta_sum_out_tmp[10][27];
        eta_sum[10][27]  = eta_sum_out_tmp[10][28];
        eta_sum[10][28]  = eta_sum_out_tmp[10][29];
        eta_sum[10][29]  = eta_sum_out_tmp[10][30];
        eta_sum[10][30]  = eta_sum_out_tmp[10][31];
        eta_sum[10][31]  = eta_sum_out_tmp[10][32];
        eta_sum[10][32]  = eta_sum_out_tmp[10][33];
        eta_sum[10][33]  = eta_sum_out_tmp[10][34];
        eta_sum[10][34]  = eta_sum_out_tmp[10][35];
        eta_sum[10][35]  = eta_sum_out_tmp[10][36];
        eta_sum[10][36]  = eta_sum_out_tmp[10][37];
        eta_sum[10][37]  = eta_sum_out_tmp[10][38];
        eta_sum[10][38]  = eta_sum_out_tmp[10][39];
        eta_sum[10][39]  = eta_sum_out_tmp[10][40];
        eta_sum[10][40]  = eta_sum_out_tmp[10][41];
    end
 
    3:begin 
        eta_sum[10][15]  = eta_sum_out_tmp[10][0];
        eta_sum[10][16]  = eta_sum_out_tmp[10][1];
        eta_sum[10][17]  = eta_sum_out_tmp[10][2];
        eta_sum[10][18]  = eta_sum_out_tmp[10][3];
        eta_sum[10][19]  = eta_sum_out_tmp[10][4];
        eta_sum[10][20]  = eta_sum_out_tmp[10][5];
        eta_sum[10][21]  = eta_sum_out_tmp[10][6];
        eta_sum[10][22]  = eta_sum_out_tmp[10][7];
        eta_sum[10][23]  = eta_sum_out_tmp[10][8];
        eta_sum[10][24]  = eta_sum_out_tmp[10][9];
        eta_sum[10][25]  = eta_sum_out_tmp[10][10];
        eta_sum[10][26]  = eta_sum_out_tmp[10][11];
        eta_sum[10][27]  = eta_sum_out_tmp[10][12];
        eta_sum[10][28]  = eta_sum_out_tmp[10][13];
        eta_sum[10][29]  = eta_sum_out_tmp[10][14];
        eta_sum[10][30]  = eta_sum_out_tmp[10][15];
        eta_sum[10][31]  = eta_sum_out_tmp[10][16];
        eta_sum[10][32]  = eta_sum_out_tmp[10][17];
        eta_sum[10][33]  = eta_sum_out_tmp[10][18];
        eta_sum[10][34]  = eta_sum_out_tmp[10][19];
        eta_sum[10][35]  = eta_sum_out_tmp[10][20];
        eta_sum[10][36]  = eta_sum_out_tmp[10][21];
        eta_sum[10][37]  = eta_sum_out_tmp[10][22];
        eta_sum[10][38]  = eta_sum_out_tmp[10][23];
        eta_sum[10][39]  = eta_sum_out_tmp[10][24];
        eta_sum[10][40]  = eta_sum_out_tmp[10][25];
        eta_sum[10][41]  = eta_sum_out_tmp[10][26];
        eta_sum[10][0]  = eta_sum_out_tmp[10][27];
        eta_sum[10][1]  = eta_sum_out_tmp[10][28];
        eta_sum[10][2]  = eta_sum_out_tmp[10][29];
        eta_sum[10][3]  = eta_sum_out_tmp[10][30];
        eta_sum[10][4]  = eta_sum_out_tmp[10][31];
        eta_sum[10][5]  = eta_sum_out_tmp[10][32];
        eta_sum[10][6]  = eta_sum_out_tmp[10][33];
        eta_sum[10][7]  = eta_sum_out_tmp[10][34];
        eta_sum[10][8]  = eta_sum_out_tmp[10][35];
        eta_sum[10][9]  = eta_sum_out_tmp[10][36];
        eta_sum[10][10]  = eta_sum_out_tmp[10][37];
        eta_sum[10][11]  = eta_sum_out_tmp[10][38];
        eta_sum[10][12]  = eta_sum_out_tmp[10][39];
        eta_sum[10][13]  = eta_sum_out_tmp[10][40];
        eta_sum[10][14]  = eta_sum_out_tmp[10][41];
    end
 
    4:begin 
        eta_sum[10][0]  = eta_sum_out_tmp[10][0];
        eta_sum[10][1]  = eta_sum_out_tmp[10][1];
        eta_sum[10][2]  = eta_sum_out_tmp[10][2];
        eta_sum[10][3]  = eta_sum_out_tmp[10][3];
        eta_sum[10][4]  = eta_sum_out_tmp[10][4];
        eta_sum[10][5]  = eta_sum_out_tmp[10][5];
        eta_sum[10][6]  = eta_sum_out_tmp[10][6];
        eta_sum[10][7]  = eta_sum_out_tmp[10][7];
        eta_sum[10][8]  = eta_sum_out_tmp[10][8];
        eta_sum[10][9]  = eta_sum_out_tmp[10][9];
        eta_sum[10][10]  = eta_sum_out_tmp[10][10];
        eta_sum[10][11]  = eta_sum_out_tmp[10][11];
        eta_sum[10][12]  = eta_sum_out_tmp[10][12];
        eta_sum[10][13]  = eta_sum_out_tmp[10][13];
        eta_sum[10][14]  = eta_sum_out_tmp[10][14];
        eta_sum[10][15]  = eta_sum_out_tmp[10][15];
        eta_sum[10][16]  = eta_sum_out_tmp[10][16];
        eta_sum[10][17]  = eta_sum_out_tmp[10][17];
        eta_sum[10][18]  = eta_sum_out_tmp[10][18];
        eta_sum[10][19]  = eta_sum_out_tmp[10][19];
        eta_sum[10][20]  = eta_sum_out_tmp[10][20];
        eta_sum[10][21]  = eta_sum_out_tmp[10][21];
        eta_sum[10][22]  = eta_sum_out_tmp[10][22];
        eta_sum[10][23]  = eta_sum_out_tmp[10][23];
        eta_sum[10][24]  = eta_sum_out_tmp[10][24];
        eta_sum[10][25]  = eta_sum_out_tmp[10][25];
        eta_sum[10][26]  = eta_sum_out_tmp[10][26];
        eta_sum[10][27]  = eta_sum_out_tmp[10][27];
        eta_sum[10][28]  = eta_sum_out_tmp[10][28];
        eta_sum[10][29]  = eta_sum_out_tmp[10][29];
        eta_sum[10][30]  = eta_sum_out_tmp[10][30];
        eta_sum[10][31]  = eta_sum_out_tmp[10][31];
        eta_sum[10][32]  = eta_sum_out_tmp[10][32];
        eta_sum[10][33]  = eta_sum_out_tmp[10][33];
        eta_sum[10][34]  = eta_sum_out_tmp[10][34];
        eta_sum[10][35]  = eta_sum_out_tmp[10][35];
        eta_sum[10][36]  = eta_sum_out_tmp[10][36];
        eta_sum[10][37]  = eta_sum_out_tmp[10][37];
        eta_sum[10][38]  = eta_sum_out_tmp[10][38];
        eta_sum[10][39]  = eta_sum_out_tmp[10][39];
        eta_sum[10][40]  = eta_sum_out_tmp[10][40];
        eta_sum[10][41]  = eta_sum_out_tmp[10][41];
    end
 
    5:begin 
        eta_sum[10][0]  = eta_sum_out_tmp[10][0];
        eta_sum[10][1]  = eta_sum_out_tmp[10][1];
        eta_sum[10][2]  = eta_sum_out_tmp[10][2];
        eta_sum[10][3]  = eta_sum_out_tmp[10][3];
        eta_sum[10][4]  = eta_sum_out_tmp[10][4];
        eta_sum[10][5]  = eta_sum_out_tmp[10][5];
        eta_sum[10][6]  = eta_sum_out_tmp[10][6];
        eta_sum[10][7]  = eta_sum_out_tmp[10][7];
        eta_sum[10][8]  = eta_sum_out_tmp[10][8];
        eta_sum[10][9]  = eta_sum_out_tmp[10][9];
        eta_sum[10][10]  = eta_sum_out_tmp[10][10];
        eta_sum[10][11]  = eta_sum_out_tmp[10][11];
        eta_sum[10][12]  = eta_sum_out_tmp[10][12];
        eta_sum[10][13]  = eta_sum_out_tmp[10][13];
        eta_sum[10][14]  = eta_sum_out_tmp[10][14];
        eta_sum[10][15]  = eta_sum_out_tmp[10][15];
        eta_sum[10][16]  = eta_sum_out_tmp[10][16];
        eta_sum[10][17]  = eta_sum_out_tmp[10][17];
        eta_sum[10][18]  = eta_sum_out_tmp[10][18];
        eta_sum[10][19]  = eta_sum_out_tmp[10][19];
        eta_sum[10][20]  = eta_sum_out_tmp[10][20];
        eta_sum[10][21]  = eta_sum_out_tmp[10][21];
        eta_sum[10][22]  = eta_sum_out_tmp[10][22];
        eta_sum[10][23]  = eta_sum_out_tmp[10][23];
        eta_sum[10][24]  = eta_sum_out_tmp[10][24];
        eta_sum[10][25]  = eta_sum_out_tmp[10][25];
        eta_sum[10][26]  = eta_sum_out_tmp[10][26];
        eta_sum[10][27]  = eta_sum_out_tmp[10][27];
        eta_sum[10][28]  = eta_sum_out_tmp[10][28];
        eta_sum[10][29]  = eta_sum_out_tmp[10][29];
        eta_sum[10][30]  = eta_sum_out_tmp[10][30];
        eta_sum[10][31]  = eta_sum_out_tmp[10][31];
        eta_sum[10][32]  = eta_sum_out_tmp[10][32];
        eta_sum[10][33]  = eta_sum_out_tmp[10][33];
        eta_sum[10][34]  = eta_sum_out_tmp[10][34];
        eta_sum[10][35]  = eta_sum_out_tmp[10][35];
        eta_sum[10][36]  = eta_sum_out_tmp[10][36];
        eta_sum[10][37]  = eta_sum_out_tmp[10][37];
        eta_sum[10][38]  = eta_sum_out_tmp[10][38];
        eta_sum[10][39]  = eta_sum_out_tmp[10][39];
        eta_sum[10][40]  = eta_sum_out_tmp[10][40];
        eta_sum[10][41]  = eta_sum_out_tmp[10][41];
    end
 
    6:begin 
        eta_sum[10][12]  = eta_sum_out_tmp[10][0];
        eta_sum[10][13]  = eta_sum_out_tmp[10][1];
        eta_sum[10][14]  = eta_sum_out_tmp[10][2];
        eta_sum[10][15]  = eta_sum_out_tmp[10][3];
        eta_sum[10][16]  = eta_sum_out_tmp[10][4];
        eta_sum[10][17]  = eta_sum_out_tmp[10][5];
        eta_sum[10][18]  = eta_sum_out_tmp[10][6];
        eta_sum[10][19]  = eta_sum_out_tmp[10][7];
        eta_sum[10][20]  = eta_sum_out_tmp[10][8];
        eta_sum[10][21]  = eta_sum_out_tmp[10][9];
        eta_sum[10][22]  = eta_sum_out_tmp[10][10];
        eta_sum[10][23]  = eta_sum_out_tmp[10][11];
        eta_sum[10][24]  = eta_sum_out_tmp[10][12];
        eta_sum[10][25]  = eta_sum_out_tmp[10][13];
        eta_sum[10][26]  = eta_sum_out_tmp[10][14];
        eta_sum[10][27]  = eta_sum_out_tmp[10][15];
        eta_sum[10][28]  = eta_sum_out_tmp[10][16];
        eta_sum[10][29]  = eta_sum_out_tmp[10][17];
        eta_sum[10][30]  = eta_sum_out_tmp[10][18];
        eta_sum[10][31]  = eta_sum_out_tmp[10][19];
        eta_sum[10][32]  = eta_sum_out_tmp[10][20];
        eta_sum[10][33]  = eta_sum_out_tmp[10][21];
        eta_sum[10][34]  = eta_sum_out_tmp[10][22];
        eta_sum[10][35]  = eta_sum_out_tmp[10][23];
        eta_sum[10][36]  = eta_sum_out_tmp[10][24];
        eta_sum[10][37]  = eta_sum_out_tmp[10][25];
        eta_sum[10][38]  = eta_sum_out_tmp[10][26];
        eta_sum[10][39]  = eta_sum_out_tmp[10][27];
        eta_sum[10][40]  = eta_sum_out_tmp[10][28];
        eta_sum[10][41]  = eta_sum_out_tmp[10][29];
        eta_sum[10][0]  = eta_sum_out_tmp[10][30];
        eta_sum[10][1]  = eta_sum_out_tmp[10][31];
        eta_sum[10][2]  = eta_sum_out_tmp[10][32];
        eta_sum[10][3]  = eta_sum_out_tmp[10][33];
        eta_sum[10][4]  = eta_sum_out_tmp[10][34];
        eta_sum[10][5]  = eta_sum_out_tmp[10][35];
        eta_sum[10][6]  = eta_sum_out_tmp[10][36];
        eta_sum[10][7]  = eta_sum_out_tmp[10][37];
        eta_sum[10][8]  = eta_sum_out_tmp[10][38];
        eta_sum[10][9]  = eta_sum_out_tmp[10][39];
        eta_sum[10][10]  = eta_sum_out_tmp[10][40];
        eta_sum[10][11]  = eta_sum_out_tmp[10][41];
    end
 
    7:begin 
        eta_sum[10][0]  = eta_sum_out_tmp[10][0];
        eta_sum[10][1]  = eta_sum_out_tmp[10][1];
        eta_sum[10][2]  = eta_sum_out_tmp[10][2];
        eta_sum[10][3]  = eta_sum_out_tmp[10][3];
        eta_sum[10][4]  = eta_sum_out_tmp[10][4];
        eta_sum[10][5]  = eta_sum_out_tmp[10][5];
        eta_sum[10][6]  = eta_sum_out_tmp[10][6];
        eta_sum[10][7]  = eta_sum_out_tmp[10][7];
        eta_sum[10][8]  = eta_sum_out_tmp[10][8];
        eta_sum[10][9]  = eta_sum_out_tmp[10][9];
        eta_sum[10][10]  = eta_sum_out_tmp[10][10];
        eta_sum[10][11]  = eta_sum_out_tmp[10][11];
        eta_sum[10][12]  = eta_sum_out_tmp[10][12];
        eta_sum[10][13]  = eta_sum_out_tmp[10][13];
        eta_sum[10][14]  = eta_sum_out_tmp[10][14];
        eta_sum[10][15]  = eta_sum_out_tmp[10][15];
        eta_sum[10][16]  = eta_sum_out_tmp[10][16];
        eta_sum[10][17]  = eta_sum_out_tmp[10][17];
        eta_sum[10][18]  = eta_sum_out_tmp[10][18];
        eta_sum[10][19]  = eta_sum_out_tmp[10][19];
        eta_sum[10][20]  = eta_sum_out_tmp[10][20];
        eta_sum[10][21]  = eta_sum_out_tmp[10][21];
        eta_sum[10][22]  = eta_sum_out_tmp[10][22];
        eta_sum[10][23]  = eta_sum_out_tmp[10][23];
        eta_sum[10][24]  = eta_sum_out_tmp[10][24];
        eta_sum[10][25]  = eta_sum_out_tmp[10][25];
        eta_sum[10][26]  = eta_sum_out_tmp[10][26];
        eta_sum[10][27]  = eta_sum_out_tmp[10][27];
        eta_sum[10][28]  = eta_sum_out_tmp[10][28];
        eta_sum[10][29]  = eta_sum_out_tmp[10][29];
        eta_sum[10][30]  = eta_sum_out_tmp[10][30];
        eta_sum[10][31]  = eta_sum_out_tmp[10][31];
        eta_sum[10][32]  = eta_sum_out_tmp[10][32];
        eta_sum[10][33]  = eta_sum_out_tmp[10][33];
        eta_sum[10][34]  = eta_sum_out_tmp[10][34];
        eta_sum[10][35]  = eta_sum_out_tmp[10][35];
        eta_sum[10][36]  = eta_sum_out_tmp[10][36];
        eta_sum[10][37]  = eta_sum_out_tmp[10][37];
        eta_sum[10][38]  = eta_sum_out_tmp[10][38];
        eta_sum[10][39]  = eta_sum_out_tmp[10][39];
        eta_sum[10][40]  = eta_sum_out_tmp[10][40];
        eta_sum[10][41]  = eta_sum_out_tmp[10][41];
    end
 
endcase
end

if (chk_n_output_valid[0] & active_cols[11]) begin
case (curr_layer)
    0:begin 
        eta_sum[11][0]  = eta_sum_out_tmp[11][0];
        eta_sum[11][1]  = eta_sum_out_tmp[11][1];
        eta_sum[11][2]  = eta_sum_out_tmp[11][2];
        eta_sum[11][3]  = eta_sum_out_tmp[11][3];
        eta_sum[11][4]  = eta_sum_out_tmp[11][4];
        eta_sum[11][5]  = eta_sum_out_tmp[11][5];
        eta_sum[11][6]  = eta_sum_out_tmp[11][6];
        eta_sum[11][7]  = eta_sum_out_tmp[11][7];
        eta_sum[11][8]  = eta_sum_out_tmp[11][8];
        eta_sum[11][9]  = eta_sum_out_tmp[11][9];
        eta_sum[11][10]  = eta_sum_out_tmp[11][10];
        eta_sum[11][11]  = eta_sum_out_tmp[11][11];
        eta_sum[11][12]  = eta_sum_out_tmp[11][12];
        eta_sum[11][13]  = eta_sum_out_tmp[11][13];
        eta_sum[11][14]  = eta_sum_out_tmp[11][14];
        eta_sum[11][15]  = eta_sum_out_tmp[11][15];
        eta_sum[11][16]  = eta_sum_out_tmp[11][16];
        eta_sum[11][17]  = eta_sum_out_tmp[11][17];
        eta_sum[11][18]  = eta_sum_out_tmp[11][18];
        eta_sum[11][19]  = eta_sum_out_tmp[11][19];
        eta_sum[11][20]  = eta_sum_out_tmp[11][20];
        eta_sum[11][21]  = eta_sum_out_tmp[11][21];
        eta_sum[11][22]  = eta_sum_out_tmp[11][22];
        eta_sum[11][23]  = eta_sum_out_tmp[11][23];
        eta_sum[11][24]  = eta_sum_out_tmp[11][24];
        eta_sum[11][25]  = eta_sum_out_tmp[11][25];
        eta_sum[11][26]  = eta_sum_out_tmp[11][26];
        eta_sum[11][27]  = eta_sum_out_tmp[11][27];
        eta_sum[11][28]  = eta_sum_out_tmp[11][28];
        eta_sum[11][29]  = eta_sum_out_tmp[11][29];
        eta_sum[11][30]  = eta_sum_out_tmp[11][30];
        eta_sum[11][31]  = eta_sum_out_tmp[11][31];
        eta_sum[11][32]  = eta_sum_out_tmp[11][32];
        eta_sum[11][33]  = eta_sum_out_tmp[11][33];
        eta_sum[11][34]  = eta_sum_out_tmp[11][34];
        eta_sum[11][35]  = eta_sum_out_tmp[11][35];
        eta_sum[11][36]  = eta_sum_out_tmp[11][36];
        eta_sum[11][37]  = eta_sum_out_tmp[11][37];
        eta_sum[11][38]  = eta_sum_out_tmp[11][38];
        eta_sum[11][39]  = eta_sum_out_tmp[11][39];
        eta_sum[11][40]  = eta_sum_out_tmp[11][40];
        eta_sum[11][41]  = eta_sum_out_tmp[11][41];
    end
 
    1:begin 
        eta_sum[11][0]  = eta_sum_out_tmp[11][0];
        eta_sum[11][1]  = eta_sum_out_tmp[11][1];
        eta_sum[11][2]  = eta_sum_out_tmp[11][2];
        eta_sum[11][3]  = eta_sum_out_tmp[11][3];
        eta_sum[11][4]  = eta_sum_out_tmp[11][4];
        eta_sum[11][5]  = eta_sum_out_tmp[11][5];
        eta_sum[11][6]  = eta_sum_out_tmp[11][6];
        eta_sum[11][7]  = eta_sum_out_tmp[11][7];
        eta_sum[11][8]  = eta_sum_out_tmp[11][8];
        eta_sum[11][9]  = eta_sum_out_tmp[11][9];
        eta_sum[11][10]  = eta_sum_out_tmp[11][10];
        eta_sum[11][11]  = eta_sum_out_tmp[11][11];
        eta_sum[11][12]  = eta_sum_out_tmp[11][12];
        eta_sum[11][13]  = eta_sum_out_tmp[11][13];
        eta_sum[11][14]  = eta_sum_out_tmp[11][14];
        eta_sum[11][15]  = eta_sum_out_tmp[11][15];
        eta_sum[11][16]  = eta_sum_out_tmp[11][16];
        eta_sum[11][17]  = eta_sum_out_tmp[11][17];
        eta_sum[11][18]  = eta_sum_out_tmp[11][18];
        eta_sum[11][19]  = eta_sum_out_tmp[11][19];
        eta_sum[11][20]  = eta_sum_out_tmp[11][20];
        eta_sum[11][21]  = eta_sum_out_tmp[11][21];
        eta_sum[11][22]  = eta_sum_out_tmp[11][22];
        eta_sum[11][23]  = eta_sum_out_tmp[11][23];
        eta_sum[11][24]  = eta_sum_out_tmp[11][24];
        eta_sum[11][25]  = eta_sum_out_tmp[11][25];
        eta_sum[11][26]  = eta_sum_out_tmp[11][26];
        eta_sum[11][27]  = eta_sum_out_tmp[11][27];
        eta_sum[11][28]  = eta_sum_out_tmp[11][28];
        eta_sum[11][29]  = eta_sum_out_tmp[11][29];
        eta_sum[11][30]  = eta_sum_out_tmp[11][30];
        eta_sum[11][31]  = eta_sum_out_tmp[11][31];
        eta_sum[11][32]  = eta_sum_out_tmp[11][32];
        eta_sum[11][33]  = eta_sum_out_tmp[11][33];
        eta_sum[11][34]  = eta_sum_out_tmp[11][34];
        eta_sum[11][35]  = eta_sum_out_tmp[11][35];
        eta_sum[11][36]  = eta_sum_out_tmp[11][36];
        eta_sum[11][37]  = eta_sum_out_tmp[11][37];
        eta_sum[11][38]  = eta_sum_out_tmp[11][38];
        eta_sum[11][39]  = eta_sum_out_tmp[11][39];
        eta_sum[11][40]  = eta_sum_out_tmp[11][40];
        eta_sum[11][41]  = eta_sum_out_tmp[11][41];
    end
 
    2:begin 
        eta_sum[11][0]  = eta_sum_out_tmp[11][0];
        eta_sum[11][1]  = eta_sum_out_tmp[11][1];
        eta_sum[11][2]  = eta_sum_out_tmp[11][2];
        eta_sum[11][3]  = eta_sum_out_tmp[11][3];
        eta_sum[11][4]  = eta_sum_out_tmp[11][4];
        eta_sum[11][5]  = eta_sum_out_tmp[11][5];
        eta_sum[11][6]  = eta_sum_out_tmp[11][6];
        eta_sum[11][7]  = eta_sum_out_tmp[11][7];
        eta_sum[11][8]  = eta_sum_out_tmp[11][8];
        eta_sum[11][9]  = eta_sum_out_tmp[11][9];
        eta_sum[11][10]  = eta_sum_out_tmp[11][10];
        eta_sum[11][11]  = eta_sum_out_tmp[11][11];
        eta_sum[11][12]  = eta_sum_out_tmp[11][12];
        eta_sum[11][13]  = eta_sum_out_tmp[11][13];
        eta_sum[11][14]  = eta_sum_out_tmp[11][14];
        eta_sum[11][15]  = eta_sum_out_tmp[11][15];
        eta_sum[11][16]  = eta_sum_out_tmp[11][16];
        eta_sum[11][17]  = eta_sum_out_tmp[11][17];
        eta_sum[11][18]  = eta_sum_out_tmp[11][18];
        eta_sum[11][19]  = eta_sum_out_tmp[11][19];
        eta_sum[11][20]  = eta_sum_out_tmp[11][20];
        eta_sum[11][21]  = eta_sum_out_tmp[11][21];
        eta_sum[11][22]  = eta_sum_out_tmp[11][22];
        eta_sum[11][23]  = eta_sum_out_tmp[11][23];
        eta_sum[11][24]  = eta_sum_out_tmp[11][24];
        eta_sum[11][25]  = eta_sum_out_tmp[11][25];
        eta_sum[11][26]  = eta_sum_out_tmp[11][26];
        eta_sum[11][27]  = eta_sum_out_tmp[11][27];
        eta_sum[11][28]  = eta_sum_out_tmp[11][28];
        eta_sum[11][29]  = eta_sum_out_tmp[11][29];
        eta_sum[11][30]  = eta_sum_out_tmp[11][30];
        eta_sum[11][31]  = eta_sum_out_tmp[11][31];
        eta_sum[11][32]  = eta_sum_out_tmp[11][32];
        eta_sum[11][33]  = eta_sum_out_tmp[11][33];
        eta_sum[11][34]  = eta_sum_out_tmp[11][34];
        eta_sum[11][35]  = eta_sum_out_tmp[11][35];
        eta_sum[11][36]  = eta_sum_out_tmp[11][36];
        eta_sum[11][37]  = eta_sum_out_tmp[11][37];
        eta_sum[11][38]  = eta_sum_out_tmp[11][38];
        eta_sum[11][39]  = eta_sum_out_tmp[11][39];
        eta_sum[11][40]  = eta_sum_out_tmp[11][40];
        eta_sum[11][41]  = eta_sum_out_tmp[11][41];
    end
 
    3:begin 
        eta_sum[11][6]  = eta_sum_out_tmp[11][0];
        eta_sum[11][7]  = eta_sum_out_tmp[11][1];
        eta_sum[11][8]  = eta_sum_out_tmp[11][2];
        eta_sum[11][9]  = eta_sum_out_tmp[11][3];
        eta_sum[11][10]  = eta_sum_out_tmp[11][4];
        eta_sum[11][11]  = eta_sum_out_tmp[11][5];
        eta_sum[11][12]  = eta_sum_out_tmp[11][6];
        eta_sum[11][13]  = eta_sum_out_tmp[11][7];
        eta_sum[11][14]  = eta_sum_out_tmp[11][8];
        eta_sum[11][15]  = eta_sum_out_tmp[11][9];
        eta_sum[11][16]  = eta_sum_out_tmp[11][10];
        eta_sum[11][17]  = eta_sum_out_tmp[11][11];
        eta_sum[11][18]  = eta_sum_out_tmp[11][12];
        eta_sum[11][19]  = eta_sum_out_tmp[11][13];
        eta_sum[11][20]  = eta_sum_out_tmp[11][14];
        eta_sum[11][21]  = eta_sum_out_tmp[11][15];
        eta_sum[11][22]  = eta_sum_out_tmp[11][16];
        eta_sum[11][23]  = eta_sum_out_tmp[11][17];
        eta_sum[11][24]  = eta_sum_out_tmp[11][18];
        eta_sum[11][25]  = eta_sum_out_tmp[11][19];
        eta_sum[11][26]  = eta_sum_out_tmp[11][20];
        eta_sum[11][27]  = eta_sum_out_tmp[11][21];
        eta_sum[11][28]  = eta_sum_out_tmp[11][22];
        eta_sum[11][29]  = eta_sum_out_tmp[11][23];
        eta_sum[11][30]  = eta_sum_out_tmp[11][24];
        eta_sum[11][31]  = eta_sum_out_tmp[11][25];
        eta_sum[11][32]  = eta_sum_out_tmp[11][26];
        eta_sum[11][33]  = eta_sum_out_tmp[11][27];
        eta_sum[11][34]  = eta_sum_out_tmp[11][28];
        eta_sum[11][35]  = eta_sum_out_tmp[11][29];
        eta_sum[11][36]  = eta_sum_out_tmp[11][30];
        eta_sum[11][37]  = eta_sum_out_tmp[11][31];
        eta_sum[11][38]  = eta_sum_out_tmp[11][32];
        eta_sum[11][39]  = eta_sum_out_tmp[11][33];
        eta_sum[11][40]  = eta_sum_out_tmp[11][34];
        eta_sum[11][41]  = eta_sum_out_tmp[11][35];
        eta_sum[11][0]  = eta_sum_out_tmp[11][36];
        eta_sum[11][1]  = eta_sum_out_tmp[11][37];
        eta_sum[11][2]  = eta_sum_out_tmp[11][38];
        eta_sum[11][3]  = eta_sum_out_tmp[11][39];
        eta_sum[11][4]  = eta_sum_out_tmp[11][40];
        eta_sum[11][5]  = eta_sum_out_tmp[11][41];
    end
 
    4:begin 
        eta_sum[11][3]  = eta_sum_out_tmp[11][0];
        eta_sum[11][4]  = eta_sum_out_tmp[11][1];
        eta_sum[11][5]  = eta_sum_out_tmp[11][2];
        eta_sum[11][6]  = eta_sum_out_tmp[11][3];
        eta_sum[11][7]  = eta_sum_out_tmp[11][4];
        eta_sum[11][8]  = eta_sum_out_tmp[11][5];
        eta_sum[11][9]  = eta_sum_out_tmp[11][6];
        eta_sum[11][10]  = eta_sum_out_tmp[11][7];
        eta_sum[11][11]  = eta_sum_out_tmp[11][8];
        eta_sum[11][12]  = eta_sum_out_tmp[11][9];
        eta_sum[11][13]  = eta_sum_out_tmp[11][10];
        eta_sum[11][14]  = eta_sum_out_tmp[11][11];
        eta_sum[11][15]  = eta_sum_out_tmp[11][12];
        eta_sum[11][16]  = eta_sum_out_tmp[11][13];
        eta_sum[11][17]  = eta_sum_out_tmp[11][14];
        eta_sum[11][18]  = eta_sum_out_tmp[11][15];
        eta_sum[11][19]  = eta_sum_out_tmp[11][16];
        eta_sum[11][20]  = eta_sum_out_tmp[11][17];
        eta_sum[11][21]  = eta_sum_out_tmp[11][18];
        eta_sum[11][22]  = eta_sum_out_tmp[11][19];
        eta_sum[11][23]  = eta_sum_out_tmp[11][20];
        eta_sum[11][24]  = eta_sum_out_tmp[11][21];
        eta_sum[11][25]  = eta_sum_out_tmp[11][22];
        eta_sum[11][26]  = eta_sum_out_tmp[11][23];
        eta_sum[11][27]  = eta_sum_out_tmp[11][24];
        eta_sum[11][28]  = eta_sum_out_tmp[11][25];
        eta_sum[11][29]  = eta_sum_out_tmp[11][26];
        eta_sum[11][30]  = eta_sum_out_tmp[11][27];
        eta_sum[11][31]  = eta_sum_out_tmp[11][28];
        eta_sum[11][32]  = eta_sum_out_tmp[11][29];
        eta_sum[11][33]  = eta_sum_out_tmp[11][30];
        eta_sum[11][34]  = eta_sum_out_tmp[11][31];
        eta_sum[11][35]  = eta_sum_out_tmp[11][32];
        eta_sum[11][36]  = eta_sum_out_tmp[11][33];
        eta_sum[11][37]  = eta_sum_out_tmp[11][34];
        eta_sum[11][38]  = eta_sum_out_tmp[11][35];
        eta_sum[11][39]  = eta_sum_out_tmp[11][36];
        eta_sum[11][40]  = eta_sum_out_tmp[11][37];
        eta_sum[11][41]  = eta_sum_out_tmp[11][38];
        eta_sum[11][0]  = eta_sum_out_tmp[11][39];
        eta_sum[11][1]  = eta_sum_out_tmp[11][40];
        eta_sum[11][2]  = eta_sum_out_tmp[11][41];
    end
 
    5:begin 
        eta_sum[11][27]  = eta_sum_out_tmp[11][0];
        eta_sum[11][28]  = eta_sum_out_tmp[11][1];
        eta_sum[11][29]  = eta_sum_out_tmp[11][2];
        eta_sum[11][30]  = eta_sum_out_tmp[11][3];
        eta_sum[11][31]  = eta_sum_out_tmp[11][4];
        eta_sum[11][32]  = eta_sum_out_tmp[11][5];
        eta_sum[11][33]  = eta_sum_out_tmp[11][6];
        eta_sum[11][34]  = eta_sum_out_tmp[11][7];
        eta_sum[11][35]  = eta_sum_out_tmp[11][8];
        eta_sum[11][36]  = eta_sum_out_tmp[11][9];
        eta_sum[11][37]  = eta_sum_out_tmp[11][10];
        eta_sum[11][38]  = eta_sum_out_tmp[11][11];
        eta_sum[11][39]  = eta_sum_out_tmp[11][12];
        eta_sum[11][40]  = eta_sum_out_tmp[11][13];
        eta_sum[11][41]  = eta_sum_out_tmp[11][14];
        eta_sum[11][0]  = eta_sum_out_tmp[11][15];
        eta_sum[11][1]  = eta_sum_out_tmp[11][16];
        eta_sum[11][2]  = eta_sum_out_tmp[11][17];
        eta_sum[11][3]  = eta_sum_out_tmp[11][18];
        eta_sum[11][4]  = eta_sum_out_tmp[11][19];
        eta_sum[11][5]  = eta_sum_out_tmp[11][20];
        eta_sum[11][6]  = eta_sum_out_tmp[11][21];
        eta_sum[11][7]  = eta_sum_out_tmp[11][22];
        eta_sum[11][8]  = eta_sum_out_tmp[11][23];
        eta_sum[11][9]  = eta_sum_out_tmp[11][24];
        eta_sum[11][10]  = eta_sum_out_tmp[11][25];
        eta_sum[11][11]  = eta_sum_out_tmp[11][26];
        eta_sum[11][12]  = eta_sum_out_tmp[11][27];
        eta_sum[11][13]  = eta_sum_out_tmp[11][28];
        eta_sum[11][14]  = eta_sum_out_tmp[11][29];
        eta_sum[11][15]  = eta_sum_out_tmp[11][30];
        eta_sum[11][16]  = eta_sum_out_tmp[11][31];
        eta_sum[11][17]  = eta_sum_out_tmp[11][32];
        eta_sum[11][18]  = eta_sum_out_tmp[11][33];
        eta_sum[11][19]  = eta_sum_out_tmp[11][34];
        eta_sum[11][20]  = eta_sum_out_tmp[11][35];
        eta_sum[11][21]  = eta_sum_out_tmp[11][36];
        eta_sum[11][22]  = eta_sum_out_tmp[11][37];
        eta_sum[11][23]  = eta_sum_out_tmp[11][38];
        eta_sum[11][24]  = eta_sum_out_tmp[11][39];
        eta_sum[11][25]  = eta_sum_out_tmp[11][40];
        eta_sum[11][26]  = eta_sum_out_tmp[11][41];
    end
 
    6:begin 
        eta_sum[11][0]  = eta_sum_out_tmp[11][0];
        eta_sum[11][1]  = eta_sum_out_tmp[11][1];
        eta_sum[11][2]  = eta_sum_out_tmp[11][2];
        eta_sum[11][3]  = eta_sum_out_tmp[11][3];
        eta_sum[11][4]  = eta_sum_out_tmp[11][4];
        eta_sum[11][5]  = eta_sum_out_tmp[11][5];
        eta_sum[11][6]  = eta_sum_out_tmp[11][6];
        eta_sum[11][7]  = eta_sum_out_tmp[11][7];
        eta_sum[11][8]  = eta_sum_out_tmp[11][8];
        eta_sum[11][9]  = eta_sum_out_tmp[11][9];
        eta_sum[11][10]  = eta_sum_out_tmp[11][10];
        eta_sum[11][11]  = eta_sum_out_tmp[11][11];
        eta_sum[11][12]  = eta_sum_out_tmp[11][12];
        eta_sum[11][13]  = eta_sum_out_tmp[11][13];
        eta_sum[11][14]  = eta_sum_out_tmp[11][14];
        eta_sum[11][15]  = eta_sum_out_tmp[11][15];
        eta_sum[11][16]  = eta_sum_out_tmp[11][16];
        eta_sum[11][17]  = eta_sum_out_tmp[11][17];
        eta_sum[11][18]  = eta_sum_out_tmp[11][18];
        eta_sum[11][19]  = eta_sum_out_tmp[11][19];
        eta_sum[11][20]  = eta_sum_out_tmp[11][20];
        eta_sum[11][21]  = eta_sum_out_tmp[11][21];
        eta_sum[11][22]  = eta_sum_out_tmp[11][22];
        eta_sum[11][23]  = eta_sum_out_tmp[11][23];
        eta_sum[11][24]  = eta_sum_out_tmp[11][24];
        eta_sum[11][25]  = eta_sum_out_tmp[11][25];
        eta_sum[11][26]  = eta_sum_out_tmp[11][26];
        eta_sum[11][27]  = eta_sum_out_tmp[11][27];
        eta_sum[11][28]  = eta_sum_out_tmp[11][28];
        eta_sum[11][29]  = eta_sum_out_tmp[11][29];
        eta_sum[11][30]  = eta_sum_out_tmp[11][30];
        eta_sum[11][31]  = eta_sum_out_tmp[11][31];
        eta_sum[11][32]  = eta_sum_out_tmp[11][32];
        eta_sum[11][33]  = eta_sum_out_tmp[11][33];
        eta_sum[11][34]  = eta_sum_out_tmp[11][34];
        eta_sum[11][35]  = eta_sum_out_tmp[11][35];
        eta_sum[11][36]  = eta_sum_out_tmp[11][36];
        eta_sum[11][37]  = eta_sum_out_tmp[11][37];
        eta_sum[11][38]  = eta_sum_out_tmp[11][38];
        eta_sum[11][39]  = eta_sum_out_tmp[11][39];
        eta_sum[11][40]  = eta_sum_out_tmp[11][40];
        eta_sum[11][41]  = eta_sum_out_tmp[11][41];
    end
 
    7:begin 
        eta_sum[11][0]  = eta_sum_out_tmp[11][0];
        eta_sum[11][1]  = eta_sum_out_tmp[11][1];
        eta_sum[11][2]  = eta_sum_out_tmp[11][2];
        eta_sum[11][3]  = eta_sum_out_tmp[11][3];
        eta_sum[11][4]  = eta_sum_out_tmp[11][4];
        eta_sum[11][5]  = eta_sum_out_tmp[11][5];
        eta_sum[11][6]  = eta_sum_out_tmp[11][6];
        eta_sum[11][7]  = eta_sum_out_tmp[11][7];
        eta_sum[11][8]  = eta_sum_out_tmp[11][8];
        eta_sum[11][9]  = eta_sum_out_tmp[11][9];
        eta_sum[11][10]  = eta_sum_out_tmp[11][10];
        eta_sum[11][11]  = eta_sum_out_tmp[11][11];
        eta_sum[11][12]  = eta_sum_out_tmp[11][12];
        eta_sum[11][13]  = eta_sum_out_tmp[11][13];
        eta_sum[11][14]  = eta_sum_out_tmp[11][14];
        eta_sum[11][15]  = eta_sum_out_tmp[11][15];
        eta_sum[11][16]  = eta_sum_out_tmp[11][16];
        eta_sum[11][17]  = eta_sum_out_tmp[11][17];
        eta_sum[11][18]  = eta_sum_out_tmp[11][18];
        eta_sum[11][19]  = eta_sum_out_tmp[11][19];
        eta_sum[11][20]  = eta_sum_out_tmp[11][20];
        eta_sum[11][21]  = eta_sum_out_tmp[11][21];
        eta_sum[11][22]  = eta_sum_out_tmp[11][22];
        eta_sum[11][23]  = eta_sum_out_tmp[11][23];
        eta_sum[11][24]  = eta_sum_out_tmp[11][24];
        eta_sum[11][25]  = eta_sum_out_tmp[11][25];
        eta_sum[11][26]  = eta_sum_out_tmp[11][26];
        eta_sum[11][27]  = eta_sum_out_tmp[11][27];
        eta_sum[11][28]  = eta_sum_out_tmp[11][28];
        eta_sum[11][29]  = eta_sum_out_tmp[11][29];
        eta_sum[11][30]  = eta_sum_out_tmp[11][30];
        eta_sum[11][31]  = eta_sum_out_tmp[11][31];
        eta_sum[11][32]  = eta_sum_out_tmp[11][32];
        eta_sum[11][33]  = eta_sum_out_tmp[11][33];
        eta_sum[11][34]  = eta_sum_out_tmp[11][34];
        eta_sum[11][35]  = eta_sum_out_tmp[11][35];
        eta_sum[11][36]  = eta_sum_out_tmp[11][36];
        eta_sum[11][37]  = eta_sum_out_tmp[11][37];
        eta_sum[11][38]  = eta_sum_out_tmp[11][38];
        eta_sum[11][39]  = eta_sum_out_tmp[11][39];
        eta_sum[11][40]  = eta_sum_out_tmp[11][40];
        eta_sum[11][41]  = eta_sum_out_tmp[11][41];
    end
 
endcase
end

if (chk_n_output_valid[0] & active_cols[12]) begin
case (curr_layer)
    0:begin 
        eta_sum[12][0]  = eta_sum_out_tmp[12][0];
        eta_sum[12][1]  = eta_sum_out_tmp[12][1];
        eta_sum[12][2]  = eta_sum_out_tmp[12][2];
        eta_sum[12][3]  = eta_sum_out_tmp[12][3];
        eta_sum[12][4]  = eta_sum_out_tmp[12][4];
        eta_sum[12][5]  = eta_sum_out_tmp[12][5];
        eta_sum[12][6]  = eta_sum_out_tmp[12][6];
        eta_sum[12][7]  = eta_sum_out_tmp[12][7];
        eta_sum[12][8]  = eta_sum_out_tmp[12][8];
        eta_sum[12][9]  = eta_sum_out_tmp[12][9];
        eta_sum[12][10]  = eta_sum_out_tmp[12][10];
        eta_sum[12][11]  = eta_sum_out_tmp[12][11];
        eta_sum[12][12]  = eta_sum_out_tmp[12][12];
        eta_sum[12][13]  = eta_sum_out_tmp[12][13];
        eta_sum[12][14]  = eta_sum_out_tmp[12][14];
        eta_sum[12][15]  = eta_sum_out_tmp[12][15];
        eta_sum[12][16]  = eta_sum_out_tmp[12][16];
        eta_sum[12][17]  = eta_sum_out_tmp[12][17];
        eta_sum[12][18]  = eta_sum_out_tmp[12][18];
        eta_sum[12][19]  = eta_sum_out_tmp[12][19];
        eta_sum[12][20]  = eta_sum_out_tmp[12][20];
        eta_sum[12][21]  = eta_sum_out_tmp[12][21];
        eta_sum[12][22]  = eta_sum_out_tmp[12][22];
        eta_sum[12][23]  = eta_sum_out_tmp[12][23];
        eta_sum[12][24]  = eta_sum_out_tmp[12][24];
        eta_sum[12][25]  = eta_sum_out_tmp[12][25];
        eta_sum[12][26]  = eta_sum_out_tmp[12][26];
        eta_sum[12][27]  = eta_sum_out_tmp[12][27];
        eta_sum[12][28]  = eta_sum_out_tmp[12][28];
        eta_sum[12][29]  = eta_sum_out_tmp[12][29];
        eta_sum[12][30]  = eta_sum_out_tmp[12][30];
        eta_sum[12][31]  = eta_sum_out_tmp[12][31];
        eta_sum[12][32]  = eta_sum_out_tmp[12][32];
        eta_sum[12][33]  = eta_sum_out_tmp[12][33];
        eta_sum[12][34]  = eta_sum_out_tmp[12][34];
        eta_sum[12][35]  = eta_sum_out_tmp[12][35];
        eta_sum[12][36]  = eta_sum_out_tmp[12][36];
        eta_sum[12][37]  = eta_sum_out_tmp[12][37];
        eta_sum[12][38]  = eta_sum_out_tmp[12][38];
        eta_sum[12][39]  = eta_sum_out_tmp[12][39];
        eta_sum[12][40]  = eta_sum_out_tmp[12][40];
        eta_sum[12][41]  = eta_sum_out_tmp[12][41];
    end
 
    1:begin 
        eta_sum[12][0]  = eta_sum_out_tmp[12][0];
        eta_sum[12][1]  = eta_sum_out_tmp[12][1];
        eta_sum[12][2]  = eta_sum_out_tmp[12][2];
        eta_sum[12][3]  = eta_sum_out_tmp[12][3];
        eta_sum[12][4]  = eta_sum_out_tmp[12][4];
        eta_sum[12][5]  = eta_sum_out_tmp[12][5];
        eta_sum[12][6]  = eta_sum_out_tmp[12][6];
        eta_sum[12][7]  = eta_sum_out_tmp[12][7];
        eta_sum[12][8]  = eta_sum_out_tmp[12][8];
        eta_sum[12][9]  = eta_sum_out_tmp[12][9];
        eta_sum[12][10]  = eta_sum_out_tmp[12][10];
        eta_sum[12][11]  = eta_sum_out_tmp[12][11];
        eta_sum[12][12]  = eta_sum_out_tmp[12][12];
        eta_sum[12][13]  = eta_sum_out_tmp[12][13];
        eta_sum[12][14]  = eta_sum_out_tmp[12][14];
        eta_sum[12][15]  = eta_sum_out_tmp[12][15];
        eta_sum[12][16]  = eta_sum_out_tmp[12][16];
        eta_sum[12][17]  = eta_sum_out_tmp[12][17];
        eta_sum[12][18]  = eta_sum_out_tmp[12][18];
        eta_sum[12][19]  = eta_sum_out_tmp[12][19];
        eta_sum[12][20]  = eta_sum_out_tmp[12][20];
        eta_sum[12][21]  = eta_sum_out_tmp[12][21];
        eta_sum[12][22]  = eta_sum_out_tmp[12][22];
        eta_sum[12][23]  = eta_sum_out_tmp[12][23];
        eta_sum[12][24]  = eta_sum_out_tmp[12][24];
        eta_sum[12][25]  = eta_sum_out_tmp[12][25];
        eta_sum[12][26]  = eta_sum_out_tmp[12][26];
        eta_sum[12][27]  = eta_sum_out_tmp[12][27];
        eta_sum[12][28]  = eta_sum_out_tmp[12][28];
        eta_sum[12][29]  = eta_sum_out_tmp[12][29];
        eta_sum[12][30]  = eta_sum_out_tmp[12][30];
        eta_sum[12][31]  = eta_sum_out_tmp[12][31];
        eta_sum[12][32]  = eta_sum_out_tmp[12][32];
        eta_sum[12][33]  = eta_sum_out_tmp[12][33];
        eta_sum[12][34]  = eta_sum_out_tmp[12][34];
        eta_sum[12][35]  = eta_sum_out_tmp[12][35];
        eta_sum[12][36]  = eta_sum_out_tmp[12][36];
        eta_sum[12][37]  = eta_sum_out_tmp[12][37];
        eta_sum[12][38]  = eta_sum_out_tmp[12][38];
        eta_sum[12][39]  = eta_sum_out_tmp[12][39];
        eta_sum[12][40]  = eta_sum_out_tmp[12][40];
        eta_sum[12][41]  = eta_sum_out_tmp[12][41];
    end
 
    2:begin 
        eta_sum[12][0]  = eta_sum_out_tmp[12][0];
        eta_sum[12][1]  = eta_sum_out_tmp[12][1];
        eta_sum[12][2]  = eta_sum_out_tmp[12][2];
        eta_sum[12][3]  = eta_sum_out_tmp[12][3];
        eta_sum[12][4]  = eta_sum_out_tmp[12][4];
        eta_sum[12][5]  = eta_sum_out_tmp[12][5];
        eta_sum[12][6]  = eta_sum_out_tmp[12][6];
        eta_sum[12][7]  = eta_sum_out_tmp[12][7];
        eta_sum[12][8]  = eta_sum_out_tmp[12][8];
        eta_sum[12][9]  = eta_sum_out_tmp[12][9];
        eta_sum[12][10]  = eta_sum_out_tmp[12][10];
        eta_sum[12][11]  = eta_sum_out_tmp[12][11];
        eta_sum[12][12]  = eta_sum_out_tmp[12][12];
        eta_sum[12][13]  = eta_sum_out_tmp[12][13];
        eta_sum[12][14]  = eta_sum_out_tmp[12][14];
        eta_sum[12][15]  = eta_sum_out_tmp[12][15];
        eta_sum[12][16]  = eta_sum_out_tmp[12][16];
        eta_sum[12][17]  = eta_sum_out_tmp[12][17];
        eta_sum[12][18]  = eta_sum_out_tmp[12][18];
        eta_sum[12][19]  = eta_sum_out_tmp[12][19];
        eta_sum[12][20]  = eta_sum_out_tmp[12][20];
        eta_sum[12][21]  = eta_sum_out_tmp[12][21];
        eta_sum[12][22]  = eta_sum_out_tmp[12][22];
        eta_sum[12][23]  = eta_sum_out_tmp[12][23];
        eta_sum[12][24]  = eta_sum_out_tmp[12][24];
        eta_sum[12][25]  = eta_sum_out_tmp[12][25];
        eta_sum[12][26]  = eta_sum_out_tmp[12][26];
        eta_sum[12][27]  = eta_sum_out_tmp[12][27];
        eta_sum[12][28]  = eta_sum_out_tmp[12][28];
        eta_sum[12][29]  = eta_sum_out_tmp[12][29];
        eta_sum[12][30]  = eta_sum_out_tmp[12][30];
        eta_sum[12][31]  = eta_sum_out_tmp[12][31];
        eta_sum[12][32]  = eta_sum_out_tmp[12][32];
        eta_sum[12][33]  = eta_sum_out_tmp[12][33];
        eta_sum[12][34]  = eta_sum_out_tmp[12][34];
        eta_sum[12][35]  = eta_sum_out_tmp[12][35];
        eta_sum[12][36]  = eta_sum_out_tmp[12][36];
        eta_sum[12][37]  = eta_sum_out_tmp[12][37];
        eta_sum[12][38]  = eta_sum_out_tmp[12][38];
        eta_sum[12][39]  = eta_sum_out_tmp[12][39];
        eta_sum[12][40]  = eta_sum_out_tmp[12][40];
        eta_sum[12][41]  = eta_sum_out_tmp[12][41];
    end
 
    3:begin 
        eta_sum[12][0]  = eta_sum_out_tmp[12][0];
        eta_sum[12][1]  = eta_sum_out_tmp[12][1];
        eta_sum[12][2]  = eta_sum_out_tmp[12][2];
        eta_sum[12][3]  = eta_sum_out_tmp[12][3];
        eta_sum[12][4]  = eta_sum_out_tmp[12][4];
        eta_sum[12][5]  = eta_sum_out_tmp[12][5];
        eta_sum[12][6]  = eta_sum_out_tmp[12][6];
        eta_sum[12][7]  = eta_sum_out_tmp[12][7];
        eta_sum[12][8]  = eta_sum_out_tmp[12][8];
        eta_sum[12][9]  = eta_sum_out_tmp[12][9];
        eta_sum[12][10]  = eta_sum_out_tmp[12][10];
        eta_sum[12][11]  = eta_sum_out_tmp[12][11];
        eta_sum[12][12]  = eta_sum_out_tmp[12][12];
        eta_sum[12][13]  = eta_sum_out_tmp[12][13];
        eta_sum[12][14]  = eta_sum_out_tmp[12][14];
        eta_sum[12][15]  = eta_sum_out_tmp[12][15];
        eta_sum[12][16]  = eta_sum_out_tmp[12][16];
        eta_sum[12][17]  = eta_sum_out_tmp[12][17];
        eta_sum[12][18]  = eta_sum_out_tmp[12][18];
        eta_sum[12][19]  = eta_sum_out_tmp[12][19];
        eta_sum[12][20]  = eta_sum_out_tmp[12][20];
        eta_sum[12][21]  = eta_sum_out_tmp[12][21];
        eta_sum[12][22]  = eta_sum_out_tmp[12][22];
        eta_sum[12][23]  = eta_sum_out_tmp[12][23];
        eta_sum[12][24]  = eta_sum_out_tmp[12][24];
        eta_sum[12][25]  = eta_sum_out_tmp[12][25];
        eta_sum[12][26]  = eta_sum_out_tmp[12][26];
        eta_sum[12][27]  = eta_sum_out_tmp[12][27];
        eta_sum[12][28]  = eta_sum_out_tmp[12][28];
        eta_sum[12][29]  = eta_sum_out_tmp[12][29];
        eta_sum[12][30]  = eta_sum_out_tmp[12][30];
        eta_sum[12][31]  = eta_sum_out_tmp[12][31];
        eta_sum[12][32]  = eta_sum_out_tmp[12][32];
        eta_sum[12][33]  = eta_sum_out_tmp[12][33];
        eta_sum[12][34]  = eta_sum_out_tmp[12][34];
        eta_sum[12][35]  = eta_sum_out_tmp[12][35];
        eta_sum[12][36]  = eta_sum_out_tmp[12][36];
        eta_sum[12][37]  = eta_sum_out_tmp[12][37];
        eta_sum[12][38]  = eta_sum_out_tmp[12][38];
        eta_sum[12][39]  = eta_sum_out_tmp[12][39];
        eta_sum[12][40]  = eta_sum_out_tmp[12][40];
        eta_sum[12][41]  = eta_sum_out_tmp[12][41];
    end
 
    4:begin 
        eta_sum[12][28]  = eta_sum_out_tmp[12][0];
        eta_sum[12][29]  = eta_sum_out_tmp[12][1];
        eta_sum[12][30]  = eta_sum_out_tmp[12][2];
        eta_sum[12][31]  = eta_sum_out_tmp[12][3];
        eta_sum[12][32]  = eta_sum_out_tmp[12][4];
        eta_sum[12][33]  = eta_sum_out_tmp[12][5];
        eta_sum[12][34]  = eta_sum_out_tmp[12][6];
        eta_sum[12][35]  = eta_sum_out_tmp[12][7];
        eta_sum[12][36]  = eta_sum_out_tmp[12][8];
        eta_sum[12][37]  = eta_sum_out_tmp[12][9];
        eta_sum[12][38]  = eta_sum_out_tmp[12][10];
        eta_sum[12][39]  = eta_sum_out_tmp[12][11];
        eta_sum[12][40]  = eta_sum_out_tmp[12][12];
        eta_sum[12][41]  = eta_sum_out_tmp[12][13];
        eta_sum[12][0]  = eta_sum_out_tmp[12][14];
        eta_sum[12][1]  = eta_sum_out_tmp[12][15];
        eta_sum[12][2]  = eta_sum_out_tmp[12][16];
        eta_sum[12][3]  = eta_sum_out_tmp[12][17];
        eta_sum[12][4]  = eta_sum_out_tmp[12][18];
        eta_sum[12][5]  = eta_sum_out_tmp[12][19];
        eta_sum[12][6]  = eta_sum_out_tmp[12][20];
        eta_sum[12][7]  = eta_sum_out_tmp[12][21];
        eta_sum[12][8]  = eta_sum_out_tmp[12][22];
        eta_sum[12][9]  = eta_sum_out_tmp[12][23];
        eta_sum[12][10]  = eta_sum_out_tmp[12][24];
        eta_sum[12][11]  = eta_sum_out_tmp[12][25];
        eta_sum[12][12]  = eta_sum_out_tmp[12][26];
        eta_sum[12][13]  = eta_sum_out_tmp[12][27];
        eta_sum[12][14]  = eta_sum_out_tmp[12][28];
        eta_sum[12][15]  = eta_sum_out_tmp[12][29];
        eta_sum[12][16]  = eta_sum_out_tmp[12][30];
        eta_sum[12][17]  = eta_sum_out_tmp[12][31];
        eta_sum[12][18]  = eta_sum_out_tmp[12][32];
        eta_sum[12][19]  = eta_sum_out_tmp[12][33];
        eta_sum[12][20]  = eta_sum_out_tmp[12][34];
        eta_sum[12][21]  = eta_sum_out_tmp[12][35];
        eta_sum[12][22]  = eta_sum_out_tmp[12][36];
        eta_sum[12][23]  = eta_sum_out_tmp[12][37];
        eta_sum[12][24]  = eta_sum_out_tmp[12][38];
        eta_sum[12][25]  = eta_sum_out_tmp[12][39];
        eta_sum[12][26]  = eta_sum_out_tmp[12][40];
        eta_sum[12][27]  = eta_sum_out_tmp[12][41];
    end
 
    5:begin 
        eta_sum[12][0]  = eta_sum_out_tmp[12][0];
        eta_sum[12][1]  = eta_sum_out_tmp[12][1];
        eta_sum[12][2]  = eta_sum_out_tmp[12][2];
        eta_sum[12][3]  = eta_sum_out_tmp[12][3];
        eta_sum[12][4]  = eta_sum_out_tmp[12][4];
        eta_sum[12][5]  = eta_sum_out_tmp[12][5];
        eta_sum[12][6]  = eta_sum_out_tmp[12][6];
        eta_sum[12][7]  = eta_sum_out_tmp[12][7];
        eta_sum[12][8]  = eta_sum_out_tmp[12][8];
        eta_sum[12][9]  = eta_sum_out_tmp[12][9];
        eta_sum[12][10]  = eta_sum_out_tmp[12][10];
        eta_sum[12][11]  = eta_sum_out_tmp[12][11];
        eta_sum[12][12]  = eta_sum_out_tmp[12][12];
        eta_sum[12][13]  = eta_sum_out_tmp[12][13];
        eta_sum[12][14]  = eta_sum_out_tmp[12][14];
        eta_sum[12][15]  = eta_sum_out_tmp[12][15];
        eta_sum[12][16]  = eta_sum_out_tmp[12][16];
        eta_sum[12][17]  = eta_sum_out_tmp[12][17];
        eta_sum[12][18]  = eta_sum_out_tmp[12][18];
        eta_sum[12][19]  = eta_sum_out_tmp[12][19];
        eta_sum[12][20]  = eta_sum_out_tmp[12][20];
        eta_sum[12][21]  = eta_sum_out_tmp[12][21];
        eta_sum[12][22]  = eta_sum_out_tmp[12][22];
        eta_sum[12][23]  = eta_sum_out_tmp[12][23];
        eta_sum[12][24]  = eta_sum_out_tmp[12][24];
        eta_sum[12][25]  = eta_sum_out_tmp[12][25];
        eta_sum[12][26]  = eta_sum_out_tmp[12][26];
        eta_sum[12][27]  = eta_sum_out_tmp[12][27];
        eta_sum[12][28]  = eta_sum_out_tmp[12][28];
        eta_sum[12][29]  = eta_sum_out_tmp[12][29];
        eta_sum[12][30]  = eta_sum_out_tmp[12][30];
        eta_sum[12][31]  = eta_sum_out_tmp[12][31];
        eta_sum[12][32]  = eta_sum_out_tmp[12][32];
        eta_sum[12][33]  = eta_sum_out_tmp[12][33];
        eta_sum[12][34]  = eta_sum_out_tmp[12][34];
        eta_sum[12][35]  = eta_sum_out_tmp[12][35];
        eta_sum[12][36]  = eta_sum_out_tmp[12][36];
        eta_sum[12][37]  = eta_sum_out_tmp[12][37];
        eta_sum[12][38]  = eta_sum_out_tmp[12][38];
        eta_sum[12][39]  = eta_sum_out_tmp[12][39];
        eta_sum[12][40]  = eta_sum_out_tmp[12][40];
        eta_sum[12][41]  = eta_sum_out_tmp[12][41];
    end
 
    6:begin 
        eta_sum[12][0]  = eta_sum_out_tmp[12][0];
        eta_sum[12][1]  = eta_sum_out_tmp[12][1];
        eta_sum[12][2]  = eta_sum_out_tmp[12][2];
        eta_sum[12][3]  = eta_sum_out_tmp[12][3];
        eta_sum[12][4]  = eta_sum_out_tmp[12][4];
        eta_sum[12][5]  = eta_sum_out_tmp[12][5];
        eta_sum[12][6]  = eta_sum_out_tmp[12][6];
        eta_sum[12][7]  = eta_sum_out_tmp[12][7];
        eta_sum[12][8]  = eta_sum_out_tmp[12][8];
        eta_sum[12][9]  = eta_sum_out_tmp[12][9];
        eta_sum[12][10]  = eta_sum_out_tmp[12][10];
        eta_sum[12][11]  = eta_sum_out_tmp[12][11];
        eta_sum[12][12]  = eta_sum_out_tmp[12][12];
        eta_sum[12][13]  = eta_sum_out_tmp[12][13];
        eta_sum[12][14]  = eta_sum_out_tmp[12][14];
        eta_sum[12][15]  = eta_sum_out_tmp[12][15];
        eta_sum[12][16]  = eta_sum_out_tmp[12][16];
        eta_sum[12][17]  = eta_sum_out_tmp[12][17];
        eta_sum[12][18]  = eta_sum_out_tmp[12][18];
        eta_sum[12][19]  = eta_sum_out_tmp[12][19];
        eta_sum[12][20]  = eta_sum_out_tmp[12][20];
        eta_sum[12][21]  = eta_sum_out_tmp[12][21];
        eta_sum[12][22]  = eta_sum_out_tmp[12][22];
        eta_sum[12][23]  = eta_sum_out_tmp[12][23];
        eta_sum[12][24]  = eta_sum_out_tmp[12][24];
        eta_sum[12][25]  = eta_sum_out_tmp[12][25];
        eta_sum[12][26]  = eta_sum_out_tmp[12][26];
        eta_sum[12][27]  = eta_sum_out_tmp[12][27];
        eta_sum[12][28]  = eta_sum_out_tmp[12][28];
        eta_sum[12][29]  = eta_sum_out_tmp[12][29];
        eta_sum[12][30]  = eta_sum_out_tmp[12][30];
        eta_sum[12][31]  = eta_sum_out_tmp[12][31];
        eta_sum[12][32]  = eta_sum_out_tmp[12][32];
        eta_sum[12][33]  = eta_sum_out_tmp[12][33];
        eta_sum[12][34]  = eta_sum_out_tmp[12][34];
        eta_sum[12][35]  = eta_sum_out_tmp[12][35];
        eta_sum[12][36]  = eta_sum_out_tmp[12][36];
        eta_sum[12][37]  = eta_sum_out_tmp[12][37];
        eta_sum[12][38]  = eta_sum_out_tmp[12][38];
        eta_sum[12][39]  = eta_sum_out_tmp[12][39];
        eta_sum[12][40]  = eta_sum_out_tmp[12][40];
        eta_sum[12][41]  = eta_sum_out_tmp[12][41];
    end
 
    7:begin 
        eta_sum[12][13]  = eta_sum_out_tmp[12][0];
        eta_sum[12][14]  = eta_sum_out_tmp[12][1];
        eta_sum[12][15]  = eta_sum_out_tmp[12][2];
        eta_sum[12][16]  = eta_sum_out_tmp[12][3];
        eta_sum[12][17]  = eta_sum_out_tmp[12][4];
        eta_sum[12][18]  = eta_sum_out_tmp[12][5];
        eta_sum[12][19]  = eta_sum_out_tmp[12][6];
        eta_sum[12][20]  = eta_sum_out_tmp[12][7];
        eta_sum[12][21]  = eta_sum_out_tmp[12][8];
        eta_sum[12][22]  = eta_sum_out_tmp[12][9];
        eta_sum[12][23]  = eta_sum_out_tmp[12][10];
        eta_sum[12][24]  = eta_sum_out_tmp[12][11];
        eta_sum[12][25]  = eta_sum_out_tmp[12][12];
        eta_sum[12][26]  = eta_sum_out_tmp[12][13];
        eta_sum[12][27]  = eta_sum_out_tmp[12][14];
        eta_sum[12][28]  = eta_sum_out_tmp[12][15];
        eta_sum[12][29]  = eta_sum_out_tmp[12][16];
        eta_sum[12][30]  = eta_sum_out_tmp[12][17];
        eta_sum[12][31]  = eta_sum_out_tmp[12][18];
        eta_sum[12][32]  = eta_sum_out_tmp[12][19];
        eta_sum[12][33]  = eta_sum_out_tmp[12][20];
        eta_sum[12][34]  = eta_sum_out_tmp[12][21];
        eta_sum[12][35]  = eta_sum_out_tmp[12][22];
        eta_sum[12][36]  = eta_sum_out_tmp[12][23];
        eta_sum[12][37]  = eta_sum_out_tmp[12][24];
        eta_sum[12][38]  = eta_sum_out_tmp[12][25];
        eta_sum[12][39]  = eta_sum_out_tmp[12][26];
        eta_sum[12][40]  = eta_sum_out_tmp[12][27];
        eta_sum[12][41]  = eta_sum_out_tmp[12][28];
        eta_sum[12][0]  = eta_sum_out_tmp[12][29];
        eta_sum[12][1]  = eta_sum_out_tmp[12][30];
        eta_sum[12][2]  = eta_sum_out_tmp[12][31];
        eta_sum[12][3]  = eta_sum_out_tmp[12][32];
        eta_sum[12][4]  = eta_sum_out_tmp[12][33];
        eta_sum[12][5]  = eta_sum_out_tmp[12][34];
        eta_sum[12][6]  = eta_sum_out_tmp[12][35];
        eta_sum[12][7]  = eta_sum_out_tmp[12][36];
        eta_sum[12][8]  = eta_sum_out_tmp[12][37];
        eta_sum[12][9]  = eta_sum_out_tmp[12][38];
        eta_sum[12][10]  = eta_sum_out_tmp[12][39];
        eta_sum[12][11]  = eta_sum_out_tmp[12][40];
        eta_sum[12][12]  = eta_sum_out_tmp[12][41];
    end
 
endcase
end

if (chk_n_output_valid[0] & active_cols[13]) begin
case (curr_layer)
    0:begin 
        eta_sum[13][0]  = eta_sum_out_tmp[13][0];
        eta_sum[13][1]  = eta_sum_out_tmp[13][1];
        eta_sum[13][2]  = eta_sum_out_tmp[13][2];
        eta_sum[13][3]  = eta_sum_out_tmp[13][3];
        eta_sum[13][4]  = eta_sum_out_tmp[13][4];
        eta_sum[13][5]  = eta_sum_out_tmp[13][5];
        eta_sum[13][6]  = eta_sum_out_tmp[13][6];
        eta_sum[13][7]  = eta_sum_out_tmp[13][7];
        eta_sum[13][8]  = eta_sum_out_tmp[13][8];
        eta_sum[13][9]  = eta_sum_out_tmp[13][9];
        eta_sum[13][10]  = eta_sum_out_tmp[13][10];
        eta_sum[13][11]  = eta_sum_out_tmp[13][11];
        eta_sum[13][12]  = eta_sum_out_tmp[13][12];
        eta_sum[13][13]  = eta_sum_out_tmp[13][13];
        eta_sum[13][14]  = eta_sum_out_tmp[13][14];
        eta_sum[13][15]  = eta_sum_out_tmp[13][15];
        eta_sum[13][16]  = eta_sum_out_tmp[13][16];
        eta_sum[13][17]  = eta_sum_out_tmp[13][17];
        eta_sum[13][18]  = eta_sum_out_tmp[13][18];
        eta_sum[13][19]  = eta_sum_out_tmp[13][19];
        eta_sum[13][20]  = eta_sum_out_tmp[13][20];
        eta_sum[13][21]  = eta_sum_out_tmp[13][21];
        eta_sum[13][22]  = eta_sum_out_tmp[13][22];
        eta_sum[13][23]  = eta_sum_out_tmp[13][23];
        eta_sum[13][24]  = eta_sum_out_tmp[13][24];
        eta_sum[13][25]  = eta_sum_out_tmp[13][25];
        eta_sum[13][26]  = eta_sum_out_tmp[13][26];
        eta_sum[13][27]  = eta_sum_out_tmp[13][27];
        eta_sum[13][28]  = eta_sum_out_tmp[13][28];
        eta_sum[13][29]  = eta_sum_out_tmp[13][29];
        eta_sum[13][30]  = eta_sum_out_tmp[13][30];
        eta_sum[13][31]  = eta_sum_out_tmp[13][31];
        eta_sum[13][32]  = eta_sum_out_tmp[13][32];
        eta_sum[13][33]  = eta_sum_out_tmp[13][33];
        eta_sum[13][34]  = eta_sum_out_tmp[13][34];
        eta_sum[13][35]  = eta_sum_out_tmp[13][35];
        eta_sum[13][36]  = eta_sum_out_tmp[13][36];
        eta_sum[13][37]  = eta_sum_out_tmp[13][37];
        eta_sum[13][38]  = eta_sum_out_tmp[13][38];
        eta_sum[13][39]  = eta_sum_out_tmp[13][39];
        eta_sum[13][40]  = eta_sum_out_tmp[13][40];
        eta_sum[13][41]  = eta_sum_out_tmp[13][41];
    end
 
    1:begin 
        eta_sum[13][0]  = eta_sum_out_tmp[13][0];
        eta_sum[13][1]  = eta_sum_out_tmp[13][1];
        eta_sum[13][2]  = eta_sum_out_tmp[13][2];
        eta_sum[13][3]  = eta_sum_out_tmp[13][3];
        eta_sum[13][4]  = eta_sum_out_tmp[13][4];
        eta_sum[13][5]  = eta_sum_out_tmp[13][5];
        eta_sum[13][6]  = eta_sum_out_tmp[13][6];
        eta_sum[13][7]  = eta_sum_out_tmp[13][7];
        eta_sum[13][8]  = eta_sum_out_tmp[13][8];
        eta_sum[13][9]  = eta_sum_out_tmp[13][9];
        eta_sum[13][10]  = eta_sum_out_tmp[13][10];
        eta_sum[13][11]  = eta_sum_out_tmp[13][11];
        eta_sum[13][12]  = eta_sum_out_tmp[13][12];
        eta_sum[13][13]  = eta_sum_out_tmp[13][13];
        eta_sum[13][14]  = eta_sum_out_tmp[13][14];
        eta_sum[13][15]  = eta_sum_out_tmp[13][15];
        eta_sum[13][16]  = eta_sum_out_tmp[13][16];
        eta_sum[13][17]  = eta_sum_out_tmp[13][17];
        eta_sum[13][18]  = eta_sum_out_tmp[13][18];
        eta_sum[13][19]  = eta_sum_out_tmp[13][19];
        eta_sum[13][20]  = eta_sum_out_tmp[13][20];
        eta_sum[13][21]  = eta_sum_out_tmp[13][21];
        eta_sum[13][22]  = eta_sum_out_tmp[13][22];
        eta_sum[13][23]  = eta_sum_out_tmp[13][23];
        eta_sum[13][24]  = eta_sum_out_tmp[13][24];
        eta_sum[13][25]  = eta_sum_out_tmp[13][25];
        eta_sum[13][26]  = eta_sum_out_tmp[13][26];
        eta_sum[13][27]  = eta_sum_out_tmp[13][27];
        eta_sum[13][28]  = eta_sum_out_tmp[13][28];
        eta_sum[13][29]  = eta_sum_out_tmp[13][29];
        eta_sum[13][30]  = eta_sum_out_tmp[13][30];
        eta_sum[13][31]  = eta_sum_out_tmp[13][31];
        eta_sum[13][32]  = eta_sum_out_tmp[13][32];
        eta_sum[13][33]  = eta_sum_out_tmp[13][33];
        eta_sum[13][34]  = eta_sum_out_tmp[13][34];
        eta_sum[13][35]  = eta_sum_out_tmp[13][35];
        eta_sum[13][36]  = eta_sum_out_tmp[13][36];
        eta_sum[13][37]  = eta_sum_out_tmp[13][37];
        eta_sum[13][38]  = eta_sum_out_tmp[13][38];
        eta_sum[13][39]  = eta_sum_out_tmp[13][39];
        eta_sum[13][40]  = eta_sum_out_tmp[13][40];
        eta_sum[13][41]  = eta_sum_out_tmp[13][41];
    end
 
    2:begin 
        eta_sum[13][0]  = eta_sum_out_tmp[13][0];
        eta_sum[13][1]  = eta_sum_out_tmp[13][1];
        eta_sum[13][2]  = eta_sum_out_tmp[13][2];
        eta_sum[13][3]  = eta_sum_out_tmp[13][3];
        eta_sum[13][4]  = eta_sum_out_tmp[13][4];
        eta_sum[13][5]  = eta_sum_out_tmp[13][5];
        eta_sum[13][6]  = eta_sum_out_tmp[13][6];
        eta_sum[13][7]  = eta_sum_out_tmp[13][7];
        eta_sum[13][8]  = eta_sum_out_tmp[13][8];
        eta_sum[13][9]  = eta_sum_out_tmp[13][9];
        eta_sum[13][10]  = eta_sum_out_tmp[13][10];
        eta_sum[13][11]  = eta_sum_out_tmp[13][11];
        eta_sum[13][12]  = eta_sum_out_tmp[13][12];
        eta_sum[13][13]  = eta_sum_out_tmp[13][13];
        eta_sum[13][14]  = eta_sum_out_tmp[13][14];
        eta_sum[13][15]  = eta_sum_out_tmp[13][15];
        eta_sum[13][16]  = eta_sum_out_tmp[13][16];
        eta_sum[13][17]  = eta_sum_out_tmp[13][17];
        eta_sum[13][18]  = eta_sum_out_tmp[13][18];
        eta_sum[13][19]  = eta_sum_out_tmp[13][19];
        eta_sum[13][20]  = eta_sum_out_tmp[13][20];
        eta_sum[13][21]  = eta_sum_out_tmp[13][21];
        eta_sum[13][22]  = eta_sum_out_tmp[13][22];
        eta_sum[13][23]  = eta_sum_out_tmp[13][23];
        eta_sum[13][24]  = eta_sum_out_tmp[13][24];
        eta_sum[13][25]  = eta_sum_out_tmp[13][25];
        eta_sum[13][26]  = eta_sum_out_tmp[13][26];
        eta_sum[13][27]  = eta_sum_out_tmp[13][27];
        eta_sum[13][28]  = eta_sum_out_tmp[13][28];
        eta_sum[13][29]  = eta_sum_out_tmp[13][29];
        eta_sum[13][30]  = eta_sum_out_tmp[13][30];
        eta_sum[13][31]  = eta_sum_out_tmp[13][31];
        eta_sum[13][32]  = eta_sum_out_tmp[13][32];
        eta_sum[13][33]  = eta_sum_out_tmp[13][33];
        eta_sum[13][34]  = eta_sum_out_tmp[13][34];
        eta_sum[13][35]  = eta_sum_out_tmp[13][35];
        eta_sum[13][36]  = eta_sum_out_tmp[13][36];
        eta_sum[13][37]  = eta_sum_out_tmp[13][37];
        eta_sum[13][38]  = eta_sum_out_tmp[13][38];
        eta_sum[13][39]  = eta_sum_out_tmp[13][39];
        eta_sum[13][40]  = eta_sum_out_tmp[13][40];
        eta_sum[13][41]  = eta_sum_out_tmp[13][41];
    end
 
    3:begin 
        eta_sum[13][0]  = eta_sum_out_tmp[13][0];
        eta_sum[13][1]  = eta_sum_out_tmp[13][1];
        eta_sum[13][2]  = eta_sum_out_tmp[13][2];
        eta_sum[13][3]  = eta_sum_out_tmp[13][3];
        eta_sum[13][4]  = eta_sum_out_tmp[13][4];
        eta_sum[13][5]  = eta_sum_out_tmp[13][5];
        eta_sum[13][6]  = eta_sum_out_tmp[13][6];
        eta_sum[13][7]  = eta_sum_out_tmp[13][7];
        eta_sum[13][8]  = eta_sum_out_tmp[13][8];
        eta_sum[13][9]  = eta_sum_out_tmp[13][9];
        eta_sum[13][10]  = eta_sum_out_tmp[13][10];
        eta_sum[13][11]  = eta_sum_out_tmp[13][11];
        eta_sum[13][12]  = eta_sum_out_tmp[13][12];
        eta_sum[13][13]  = eta_sum_out_tmp[13][13];
        eta_sum[13][14]  = eta_sum_out_tmp[13][14];
        eta_sum[13][15]  = eta_sum_out_tmp[13][15];
        eta_sum[13][16]  = eta_sum_out_tmp[13][16];
        eta_sum[13][17]  = eta_sum_out_tmp[13][17];
        eta_sum[13][18]  = eta_sum_out_tmp[13][18];
        eta_sum[13][19]  = eta_sum_out_tmp[13][19];
        eta_sum[13][20]  = eta_sum_out_tmp[13][20];
        eta_sum[13][21]  = eta_sum_out_tmp[13][21];
        eta_sum[13][22]  = eta_sum_out_tmp[13][22];
        eta_sum[13][23]  = eta_sum_out_tmp[13][23];
        eta_sum[13][24]  = eta_sum_out_tmp[13][24];
        eta_sum[13][25]  = eta_sum_out_tmp[13][25];
        eta_sum[13][26]  = eta_sum_out_tmp[13][26];
        eta_sum[13][27]  = eta_sum_out_tmp[13][27];
        eta_sum[13][28]  = eta_sum_out_tmp[13][28];
        eta_sum[13][29]  = eta_sum_out_tmp[13][29];
        eta_sum[13][30]  = eta_sum_out_tmp[13][30];
        eta_sum[13][31]  = eta_sum_out_tmp[13][31];
        eta_sum[13][32]  = eta_sum_out_tmp[13][32];
        eta_sum[13][33]  = eta_sum_out_tmp[13][33];
        eta_sum[13][34]  = eta_sum_out_tmp[13][34];
        eta_sum[13][35]  = eta_sum_out_tmp[13][35];
        eta_sum[13][36]  = eta_sum_out_tmp[13][36];
        eta_sum[13][37]  = eta_sum_out_tmp[13][37];
        eta_sum[13][38]  = eta_sum_out_tmp[13][38];
        eta_sum[13][39]  = eta_sum_out_tmp[13][39];
        eta_sum[13][40]  = eta_sum_out_tmp[13][40];
        eta_sum[13][41]  = eta_sum_out_tmp[13][41];
    end
 
    4:begin 
        eta_sum[13][0]  = eta_sum_out_tmp[13][0];
        eta_sum[13][1]  = eta_sum_out_tmp[13][1];
        eta_sum[13][2]  = eta_sum_out_tmp[13][2];
        eta_sum[13][3]  = eta_sum_out_tmp[13][3];
        eta_sum[13][4]  = eta_sum_out_tmp[13][4];
        eta_sum[13][5]  = eta_sum_out_tmp[13][5];
        eta_sum[13][6]  = eta_sum_out_tmp[13][6];
        eta_sum[13][7]  = eta_sum_out_tmp[13][7];
        eta_sum[13][8]  = eta_sum_out_tmp[13][8];
        eta_sum[13][9]  = eta_sum_out_tmp[13][9];
        eta_sum[13][10]  = eta_sum_out_tmp[13][10];
        eta_sum[13][11]  = eta_sum_out_tmp[13][11];
        eta_sum[13][12]  = eta_sum_out_tmp[13][12];
        eta_sum[13][13]  = eta_sum_out_tmp[13][13];
        eta_sum[13][14]  = eta_sum_out_tmp[13][14];
        eta_sum[13][15]  = eta_sum_out_tmp[13][15];
        eta_sum[13][16]  = eta_sum_out_tmp[13][16];
        eta_sum[13][17]  = eta_sum_out_tmp[13][17];
        eta_sum[13][18]  = eta_sum_out_tmp[13][18];
        eta_sum[13][19]  = eta_sum_out_tmp[13][19];
        eta_sum[13][20]  = eta_sum_out_tmp[13][20];
        eta_sum[13][21]  = eta_sum_out_tmp[13][21];
        eta_sum[13][22]  = eta_sum_out_tmp[13][22];
        eta_sum[13][23]  = eta_sum_out_tmp[13][23];
        eta_sum[13][24]  = eta_sum_out_tmp[13][24];
        eta_sum[13][25]  = eta_sum_out_tmp[13][25];
        eta_sum[13][26]  = eta_sum_out_tmp[13][26];
        eta_sum[13][27]  = eta_sum_out_tmp[13][27];
        eta_sum[13][28]  = eta_sum_out_tmp[13][28];
        eta_sum[13][29]  = eta_sum_out_tmp[13][29];
        eta_sum[13][30]  = eta_sum_out_tmp[13][30];
        eta_sum[13][31]  = eta_sum_out_tmp[13][31];
        eta_sum[13][32]  = eta_sum_out_tmp[13][32];
        eta_sum[13][33]  = eta_sum_out_tmp[13][33];
        eta_sum[13][34]  = eta_sum_out_tmp[13][34];
        eta_sum[13][35]  = eta_sum_out_tmp[13][35];
        eta_sum[13][36]  = eta_sum_out_tmp[13][36];
        eta_sum[13][37]  = eta_sum_out_tmp[13][37];
        eta_sum[13][38]  = eta_sum_out_tmp[13][38];
        eta_sum[13][39]  = eta_sum_out_tmp[13][39];
        eta_sum[13][40]  = eta_sum_out_tmp[13][40];
        eta_sum[13][41]  = eta_sum_out_tmp[13][41];
    end
 
    5:begin 
        eta_sum[13][23]  = eta_sum_out_tmp[13][0];
        eta_sum[13][24]  = eta_sum_out_tmp[13][1];
        eta_sum[13][25]  = eta_sum_out_tmp[13][2];
        eta_sum[13][26]  = eta_sum_out_tmp[13][3];
        eta_sum[13][27]  = eta_sum_out_tmp[13][4];
        eta_sum[13][28]  = eta_sum_out_tmp[13][5];
        eta_sum[13][29]  = eta_sum_out_tmp[13][6];
        eta_sum[13][30]  = eta_sum_out_tmp[13][7];
        eta_sum[13][31]  = eta_sum_out_tmp[13][8];
        eta_sum[13][32]  = eta_sum_out_tmp[13][9];
        eta_sum[13][33]  = eta_sum_out_tmp[13][10];
        eta_sum[13][34]  = eta_sum_out_tmp[13][11];
        eta_sum[13][35]  = eta_sum_out_tmp[13][12];
        eta_sum[13][36]  = eta_sum_out_tmp[13][13];
        eta_sum[13][37]  = eta_sum_out_tmp[13][14];
        eta_sum[13][38]  = eta_sum_out_tmp[13][15];
        eta_sum[13][39]  = eta_sum_out_tmp[13][16];
        eta_sum[13][40]  = eta_sum_out_tmp[13][17];
        eta_sum[13][41]  = eta_sum_out_tmp[13][18];
        eta_sum[13][0]  = eta_sum_out_tmp[13][19];
        eta_sum[13][1]  = eta_sum_out_tmp[13][20];
        eta_sum[13][2]  = eta_sum_out_tmp[13][21];
        eta_sum[13][3]  = eta_sum_out_tmp[13][22];
        eta_sum[13][4]  = eta_sum_out_tmp[13][23];
        eta_sum[13][5]  = eta_sum_out_tmp[13][24];
        eta_sum[13][6]  = eta_sum_out_tmp[13][25];
        eta_sum[13][7]  = eta_sum_out_tmp[13][26];
        eta_sum[13][8]  = eta_sum_out_tmp[13][27];
        eta_sum[13][9]  = eta_sum_out_tmp[13][28];
        eta_sum[13][10]  = eta_sum_out_tmp[13][29];
        eta_sum[13][11]  = eta_sum_out_tmp[13][30];
        eta_sum[13][12]  = eta_sum_out_tmp[13][31];
        eta_sum[13][13]  = eta_sum_out_tmp[13][32];
        eta_sum[13][14]  = eta_sum_out_tmp[13][33];
        eta_sum[13][15]  = eta_sum_out_tmp[13][34];
        eta_sum[13][16]  = eta_sum_out_tmp[13][35];
        eta_sum[13][17]  = eta_sum_out_tmp[13][36];
        eta_sum[13][18]  = eta_sum_out_tmp[13][37];
        eta_sum[13][19]  = eta_sum_out_tmp[13][38];
        eta_sum[13][20]  = eta_sum_out_tmp[13][39];
        eta_sum[13][21]  = eta_sum_out_tmp[13][40];
        eta_sum[13][22]  = eta_sum_out_tmp[13][41];
    end
 
    6:begin 
        eta_sum[13][0]  = eta_sum_out_tmp[13][0];
        eta_sum[13][1]  = eta_sum_out_tmp[13][1];
        eta_sum[13][2]  = eta_sum_out_tmp[13][2];
        eta_sum[13][3]  = eta_sum_out_tmp[13][3];
        eta_sum[13][4]  = eta_sum_out_tmp[13][4];
        eta_sum[13][5]  = eta_sum_out_tmp[13][5];
        eta_sum[13][6]  = eta_sum_out_tmp[13][6];
        eta_sum[13][7]  = eta_sum_out_tmp[13][7];
        eta_sum[13][8]  = eta_sum_out_tmp[13][8];
        eta_sum[13][9]  = eta_sum_out_tmp[13][9];
        eta_sum[13][10]  = eta_sum_out_tmp[13][10];
        eta_sum[13][11]  = eta_sum_out_tmp[13][11];
        eta_sum[13][12]  = eta_sum_out_tmp[13][12];
        eta_sum[13][13]  = eta_sum_out_tmp[13][13];
        eta_sum[13][14]  = eta_sum_out_tmp[13][14];
        eta_sum[13][15]  = eta_sum_out_tmp[13][15];
        eta_sum[13][16]  = eta_sum_out_tmp[13][16];
        eta_sum[13][17]  = eta_sum_out_tmp[13][17];
        eta_sum[13][18]  = eta_sum_out_tmp[13][18];
        eta_sum[13][19]  = eta_sum_out_tmp[13][19];
        eta_sum[13][20]  = eta_sum_out_tmp[13][20];
        eta_sum[13][21]  = eta_sum_out_tmp[13][21];
        eta_sum[13][22]  = eta_sum_out_tmp[13][22];
        eta_sum[13][23]  = eta_sum_out_tmp[13][23];
        eta_sum[13][24]  = eta_sum_out_tmp[13][24];
        eta_sum[13][25]  = eta_sum_out_tmp[13][25];
        eta_sum[13][26]  = eta_sum_out_tmp[13][26];
        eta_sum[13][27]  = eta_sum_out_tmp[13][27];
        eta_sum[13][28]  = eta_sum_out_tmp[13][28];
        eta_sum[13][29]  = eta_sum_out_tmp[13][29];
        eta_sum[13][30]  = eta_sum_out_tmp[13][30];
        eta_sum[13][31]  = eta_sum_out_tmp[13][31];
        eta_sum[13][32]  = eta_sum_out_tmp[13][32];
        eta_sum[13][33]  = eta_sum_out_tmp[13][33];
        eta_sum[13][34]  = eta_sum_out_tmp[13][34];
        eta_sum[13][35]  = eta_sum_out_tmp[13][35];
        eta_sum[13][36]  = eta_sum_out_tmp[13][36];
        eta_sum[13][37]  = eta_sum_out_tmp[13][37];
        eta_sum[13][38]  = eta_sum_out_tmp[13][38];
        eta_sum[13][39]  = eta_sum_out_tmp[13][39];
        eta_sum[13][40]  = eta_sum_out_tmp[13][40];
        eta_sum[13][41]  = eta_sum_out_tmp[13][41];
    end
 
    7:begin 
        eta_sum[13][0]  = eta_sum_out_tmp[13][0];
        eta_sum[13][1]  = eta_sum_out_tmp[13][1];
        eta_sum[13][2]  = eta_sum_out_tmp[13][2];
        eta_sum[13][3]  = eta_sum_out_tmp[13][3];
        eta_sum[13][4]  = eta_sum_out_tmp[13][4];
        eta_sum[13][5]  = eta_sum_out_tmp[13][5];
        eta_sum[13][6]  = eta_sum_out_tmp[13][6];
        eta_sum[13][7]  = eta_sum_out_tmp[13][7];
        eta_sum[13][8]  = eta_sum_out_tmp[13][8];
        eta_sum[13][9]  = eta_sum_out_tmp[13][9];
        eta_sum[13][10]  = eta_sum_out_tmp[13][10];
        eta_sum[13][11]  = eta_sum_out_tmp[13][11];
        eta_sum[13][12]  = eta_sum_out_tmp[13][12];
        eta_sum[13][13]  = eta_sum_out_tmp[13][13];
        eta_sum[13][14]  = eta_sum_out_tmp[13][14];
        eta_sum[13][15]  = eta_sum_out_tmp[13][15];
        eta_sum[13][16]  = eta_sum_out_tmp[13][16];
        eta_sum[13][17]  = eta_sum_out_tmp[13][17];
        eta_sum[13][18]  = eta_sum_out_tmp[13][18];
        eta_sum[13][19]  = eta_sum_out_tmp[13][19];
        eta_sum[13][20]  = eta_sum_out_tmp[13][20];
        eta_sum[13][21]  = eta_sum_out_tmp[13][21];
        eta_sum[13][22]  = eta_sum_out_tmp[13][22];
        eta_sum[13][23]  = eta_sum_out_tmp[13][23];
        eta_sum[13][24]  = eta_sum_out_tmp[13][24];
        eta_sum[13][25]  = eta_sum_out_tmp[13][25];
        eta_sum[13][26]  = eta_sum_out_tmp[13][26];
        eta_sum[13][27]  = eta_sum_out_tmp[13][27];
        eta_sum[13][28]  = eta_sum_out_tmp[13][28];
        eta_sum[13][29]  = eta_sum_out_tmp[13][29];
        eta_sum[13][30]  = eta_sum_out_tmp[13][30];
        eta_sum[13][31]  = eta_sum_out_tmp[13][31];
        eta_sum[13][32]  = eta_sum_out_tmp[13][32];
        eta_sum[13][33]  = eta_sum_out_tmp[13][33];
        eta_sum[13][34]  = eta_sum_out_tmp[13][34];
        eta_sum[13][35]  = eta_sum_out_tmp[13][35];
        eta_sum[13][36]  = eta_sum_out_tmp[13][36];
        eta_sum[13][37]  = eta_sum_out_tmp[13][37];
        eta_sum[13][38]  = eta_sum_out_tmp[13][38];
        eta_sum[13][39]  = eta_sum_out_tmp[13][39];
        eta_sum[13][40]  = eta_sum_out_tmp[13][40];
        eta_sum[13][41]  = eta_sum_out_tmp[13][41];
    end
 
endcase
end

if (chk_n_output_valid[0] & active_cols[14]) begin
case (curr_layer)
    0:begin 
        eta_sum[14][0]  = eta_sum_out_tmp[14][0];
        eta_sum[14][1]  = eta_sum_out_tmp[14][1];
        eta_sum[14][2]  = eta_sum_out_tmp[14][2];
        eta_sum[14][3]  = eta_sum_out_tmp[14][3];
        eta_sum[14][4]  = eta_sum_out_tmp[14][4];
        eta_sum[14][5]  = eta_sum_out_tmp[14][5];
        eta_sum[14][6]  = eta_sum_out_tmp[14][6];
        eta_sum[14][7]  = eta_sum_out_tmp[14][7];
        eta_sum[14][8]  = eta_sum_out_tmp[14][8];
        eta_sum[14][9]  = eta_sum_out_tmp[14][9];
        eta_sum[14][10]  = eta_sum_out_tmp[14][10];
        eta_sum[14][11]  = eta_sum_out_tmp[14][11];
        eta_sum[14][12]  = eta_sum_out_tmp[14][12];
        eta_sum[14][13]  = eta_sum_out_tmp[14][13];
        eta_sum[14][14]  = eta_sum_out_tmp[14][14];
        eta_sum[14][15]  = eta_sum_out_tmp[14][15];
        eta_sum[14][16]  = eta_sum_out_tmp[14][16];
        eta_sum[14][17]  = eta_sum_out_tmp[14][17];
        eta_sum[14][18]  = eta_sum_out_tmp[14][18];
        eta_sum[14][19]  = eta_sum_out_tmp[14][19];
        eta_sum[14][20]  = eta_sum_out_tmp[14][20];
        eta_sum[14][21]  = eta_sum_out_tmp[14][21];
        eta_sum[14][22]  = eta_sum_out_tmp[14][22];
        eta_sum[14][23]  = eta_sum_out_tmp[14][23];
        eta_sum[14][24]  = eta_sum_out_tmp[14][24];
        eta_sum[14][25]  = eta_sum_out_tmp[14][25];
        eta_sum[14][26]  = eta_sum_out_tmp[14][26];
        eta_sum[14][27]  = eta_sum_out_tmp[14][27];
        eta_sum[14][28]  = eta_sum_out_tmp[14][28];
        eta_sum[14][29]  = eta_sum_out_tmp[14][29];
        eta_sum[14][30]  = eta_sum_out_tmp[14][30];
        eta_sum[14][31]  = eta_sum_out_tmp[14][31];
        eta_sum[14][32]  = eta_sum_out_tmp[14][32];
        eta_sum[14][33]  = eta_sum_out_tmp[14][33];
        eta_sum[14][34]  = eta_sum_out_tmp[14][34];
        eta_sum[14][35]  = eta_sum_out_tmp[14][35];
        eta_sum[14][36]  = eta_sum_out_tmp[14][36];
        eta_sum[14][37]  = eta_sum_out_tmp[14][37];
        eta_sum[14][38]  = eta_sum_out_tmp[14][38];
        eta_sum[14][39]  = eta_sum_out_tmp[14][39];
        eta_sum[14][40]  = eta_sum_out_tmp[14][40];
        eta_sum[14][41]  = eta_sum_out_tmp[14][41];
    end
 
    1:begin 
        eta_sum[14][0]  = eta_sum_out_tmp[14][0];
        eta_sum[14][1]  = eta_sum_out_tmp[14][1];
        eta_sum[14][2]  = eta_sum_out_tmp[14][2];
        eta_sum[14][3]  = eta_sum_out_tmp[14][3];
        eta_sum[14][4]  = eta_sum_out_tmp[14][4];
        eta_sum[14][5]  = eta_sum_out_tmp[14][5];
        eta_sum[14][6]  = eta_sum_out_tmp[14][6];
        eta_sum[14][7]  = eta_sum_out_tmp[14][7];
        eta_sum[14][8]  = eta_sum_out_tmp[14][8];
        eta_sum[14][9]  = eta_sum_out_tmp[14][9];
        eta_sum[14][10]  = eta_sum_out_tmp[14][10];
        eta_sum[14][11]  = eta_sum_out_tmp[14][11];
        eta_sum[14][12]  = eta_sum_out_tmp[14][12];
        eta_sum[14][13]  = eta_sum_out_tmp[14][13];
        eta_sum[14][14]  = eta_sum_out_tmp[14][14];
        eta_sum[14][15]  = eta_sum_out_tmp[14][15];
        eta_sum[14][16]  = eta_sum_out_tmp[14][16];
        eta_sum[14][17]  = eta_sum_out_tmp[14][17];
        eta_sum[14][18]  = eta_sum_out_tmp[14][18];
        eta_sum[14][19]  = eta_sum_out_tmp[14][19];
        eta_sum[14][20]  = eta_sum_out_tmp[14][20];
        eta_sum[14][21]  = eta_sum_out_tmp[14][21];
        eta_sum[14][22]  = eta_sum_out_tmp[14][22];
        eta_sum[14][23]  = eta_sum_out_tmp[14][23];
        eta_sum[14][24]  = eta_sum_out_tmp[14][24];
        eta_sum[14][25]  = eta_sum_out_tmp[14][25];
        eta_sum[14][26]  = eta_sum_out_tmp[14][26];
        eta_sum[14][27]  = eta_sum_out_tmp[14][27];
        eta_sum[14][28]  = eta_sum_out_tmp[14][28];
        eta_sum[14][29]  = eta_sum_out_tmp[14][29];
        eta_sum[14][30]  = eta_sum_out_tmp[14][30];
        eta_sum[14][31]  = eta_sum_out_tmp[14][31];
        eta_sum[14][32]  = eta_sum_out_tmp[14][32];
        eta_sum[14][33]  = eta_sum_out_tmp[14][33];
        eta_sum[14][34]  = eta_sum_out_tmp[14][34];
        eta_sum[14][35]  = eta_sum_out_tmp[14][35];
        eta_sum[14][36]  = eta_sum_out_tmp[14][36];
        eta_sum[14][37]  = eta_sum_out_tmp[14][37];
        eta_sum[14][38]  = eta_sum_out_tmp[14][38];
        eta_sum[14][39]  = eta_sum_out_tmp[14][39];
        eta_sum[14][40]  = eta_sum_out_tmp[14][40];
        eta_sum[14][41]  = eta_sum_out_tmp[14][41];
    end
 
    2:begin 
        eta_sum[14][0]  = eta_sum_out_tmp[14][0];
        eta_sum[14][1]  = eta_sum_out_tmp[14][1];
        eta_sum[14][2]  = eta_sum_out_tmp[14][2];
        eta_sum[14][3]  = eta_sum_out_tmp[14][3];
        eta_sum[14][4]  = eta_sum_out_tmp[14][4];
        eta_sum[14][5]  = eta_sum_out_tmp[14][5];
        eta_sum[14][6]  = eta_sum_out_tmp[14][6];
        eta_sum[14][7]  = eta_sum_out_tmp[14][7];
        eta_sum[14][8]  = eta_sum_out_tmp[14][8];
        eta_sum[14][9]  = eta_sum_out_tmp[14][9];
        eta_sum[14][10]  = eta_sum_out_tmp[14][10];
        eta_sum[14][11]  = eta_sum_out_tmp[14][11];
        eta_sum[14][12]  = eta_sum_out_tmp[14][12];
        eta_sum[14][13]  = eta_sum_out_tmp[14][13];
        eta_sum[14][14]  = eta_sum_out_tmp[14][14];
        eta_sum[14][15]  = eta_sum_out_tmp[14][15];
        eta_sum[14][16]  = eta_sum_out_tmp[14][16];
        eta_sum[14][17]  = eta_sum_out_tmp[14][17];
        eta_sum[14][18]  = eta_sum_out_tmp[14][18];
        eta_sum[14][19]  = eta_sum_out_tmp[14][19];
        eta_sum[14][20]  = eta_sum_out_tmp[14][20];
        eta_sum[14][21]  = eta_sum_out_tmp[14][21];
        eta_sum[14][22]  = eta_sum_out_tmp[14][22];
        eta_sum[14][23]  = eta_sum_out_tmp[14][23];
        eta_sum[14][24]  = eta_sum_out_tmp[14][24];
        eta_sum[14][25]  = eta_sum_out_tmp[14][25];
        eta_sum[14][26]  = eta_sum_out_tmp[14][26];
        eta_sum[14][27]  = eta_sum_out_tmp[14][27];
        eta_sum[14][28]  = eta_sum_out_tmp[14][28];
        eta_sum[14][29]  = eta_sum_out_tmp[14][29];
        eta_sum[14][30]  = eta_sum_out_tmp[14][30];
        eta_sum[14][31]  = eta_sum_out_tmp[14][31];
        eta_sum[14][32]  = eta_sum_out_tmp[14][32];
        eta_sum[14][33]  = eta_sum_out_tmp[14][33];
        eta_sum[14][34]  = eta_sum_out_tmp[14][34];
        eta_sum[14][35]  = eta_sum_out_tmp[14][35];
        eta_sum[14][36]  = eta_sum_out_tmp[14][36];
        eta_sum[14][37]  = eta_sum_out_tmp[14][37];
        eta_sum[14][38]  = eta_sum_out_tmp[14][38];
        eta_sum[14][39]  = eta_sum_out_tmp[14][39];
        eta_sum[14][40]  = eta_sum_out_tmp[14][40];
        eta_sum[14][41]  = eta_sum_out_tmp[14][41];
    end
 
    3:begin 
        eta_sum[14][0]  = eta_sum_out_tmp[14][0];
        eta_sum[14][1]  = eta_sum_out_tmp[14][1];
        eta_sum[14][2]  = eta_sum_out_tmp[14][2];
        eta_sum[14][3]  = eta_sum_out_tmp[14][3];
        eta_sum[14][4]  = eta_sum_out_tmp[14][4];
        eta_sum[14][5]  = eta_sum_out_tmp[14][5];
        eta_sum[14][6]  = eta_sum_out_tmp[14][6];
        eta_sum[14][7]  = eta_sum_out_tmp[14][7];
        eta_sum[14][8]  = eta_sum_out_tmp[14][8];
        eta_sum[14][9]  = eta_sum_out_tmp[14][9];
        eta_sum[14][10]  = eta_sum_out_tmp[14][10];
        eta_sum[14][11]  = eta_sum_out_tmp[14][11];
        eta_sum[14][12]  = eta_sum_out_tmp[14][12];
        eta_sum[14][13]  = eta_sum_out_tmp[14][13];
        eta_sum[14][14]  = eta_sum_out_tmp[14][14];
        eta_sum[14][15]  = eta_sum_out_tmp[14][15];
        eta_sum[14][16]  = eta_sum_out_tmp[14][16];
        eta_sum[14][17]  = eta_sum_out_tmp[14][17];
        eta_sum[14][18]  = eta_sum_out_tmp[14][18];
        eta_sum[14][19]  = eta_sum_out_tmp[14][19];
        eta_sum[14][20]  = eta_sum_out_tmp[14][20];
        eta_sum[14][21]  = eta_sum_out_tmp[14][21];
        eta_sum[14][22]  = eta_sum_out_tmp[14][22];
        eta_sum[14][23]  = eta_sum_out_tmp[14][23];
        eta_sum[14][24]  = eta_sum_out_tmp[14][24];
        eta_sum[14][25]  = eta_sum_out_tmp[14][25];
        eta_sum[14][26]  = eta_sum_out_tmp[14][26];
        eta_sum[14][27]  = eta_sum_out_tmp[14][27];
        eta_sum[14][28]  = eta_sum_out_tmp[14][28];
        eta_sum[14][29]  = eta_sum_out_tmp[14][29];
        eta_sum[14][30]  = eta_sum_out_tmp[14][30];
        eta_sum[14][31]  = eta_sum_out_tmp[14][31];
        eta_sum[14][32]  = eta_sum_out_tmp[14][32];
        eta_sum[14][33]  = eta_sum_out_tmp[14][33];
        eta_sum[14][34]  = eta_sum_out_tmp[14][34];
        eta_sum[14][35]  = eta_sum_out_tmp[14][35];
        eta_sum[14][36]  = eta_sum_out_tmp[14][36];
        eta_sum[14][37]  = eta_sum_out_tmp[14][37];
        eta_sum[14][38]  = eta_sum_out_tmp[14][38];
        eta_sum[14][39]  = eta_sum_out_tmp[14][39];
        eta_sum[14][40]  = eta_sum_out_tmp[14][40];
        eta_sum[14][41]  = eta_sum_out_tmp[14][41];
    end
 
    4:begin 
        eta_sum[14][0]  = eta_sum_out_tmp[14][0];
        eta_sum[14][1]  = eta_sum_out_tmp[14][1];
        eta_sum[14][2]  = eta_sum_out_tmp[14][2];
        eta_sum[14][3]  = eta_sum_out_tmp[14][3];
        eta_sum[14][4]  = eta_sum_out_tmp[14][4];
        eta_sum[14][5]  = eta_sum_out_tmp[14][5];
        eta_sum[14][6]  = eta_sum_out_tmp[14][6];
        eta_sum[14][7]  = eta_sum_out_tmp[14][7];
        eta_sum[14][8]  = eta_sum_out_tmp[14][8];
        eta_sum[14][9]  = eta_sum_out_tmp[14][9];
        eta_sum[14][10]  = eta_sum_out_tmp[14][10];
        eta_sum[14][11]  = eta_sum_out_tmp[14][11];
        eta_sum[14][12]  = eta_sum_out_tmp[14][12];
        eta_sum[14][13]  = eta_sum_out_tmp[14][13];
        eta_sum[14][14]  = eta_sum_out_tmp[14][14];
        eta_sum[14][15]  = eta_sum_out_tmp[14][15];
        eta_sum[14][16]  = eta_sum_out_tmp[14][16];
        eta_sum[14][17]  = eta_sum_out_tmp[14][17];
        eta_sum[14][18]  = eta_sum_out_tmp[14][18];
        eta_sum[14][19]  = eta_sum_out_tmp[14][19];
        eta_sum[14][20]  = eta_sum_out_tmp[14][20];
        eta_sum[14][21]  = eta_sum_out_tmp[14][21];
        eta_sum[14][22]  = eta_sum_out_tmp[14][22];
        eta_sum[14][23]  = eta_sum_out_tmp[14][23];
        eta_sum[14][24]  = eta_sum_out_tmp[14][24];
        eta_sum[14][25]  = eta_sum_out_tmp[14][25];
        eta_sum[14][26]  = eta_sum_out_tmp[14][26];
        eta_sum[14][27]  = eta_sum_out_tmp[14][27];
        eta_sum[14][28]  = eta_sum_out_tmp[14][28];
        eta_sum[14][29]  = eta_sum_out_tmp[14][29];
        eta_sum[14][30]  = eta_sum_out_tmp[14][30];
        eta_sum[14][31]  = eta_sum_out_tmp[14][31];
        eta_sum[14][32]  = eta_sum_out_tmp[14][32];
        eta_sum[14][33]  = eta_sum_out_tmp[14][33];
        eta_sum[14][34]  = eta_sum_out_tmp[14][34];
        eta_sum[14][35]  = eta_sum_out_tmp[14][35];
        eta_sum[14][36]  = eta_sum_out_tmp[14][36];
        eta_sum[14][37]  = eta_sum_out_tmp[14][37];
        eta_sum[14][38]  = eta_sum_out_tmp[14][38];
        eta_sum[14][39]  = eta_sum_out_tmp[14][39];
        eta_sum[14][40]  = eta_sum_out_tmp[14][40];
        eta_sum[14][41]  = eta_sum_out_tmp[14][41];
    end
 
    5:begin 
        eta_sum[14][0]  = eta_sum_out_tmp[14][0];
        eta_sum[14][1]  = eta_sum_out_tmp[14][1];
        eta_sum[14][2]  = eta_sum_out_tmp[14][2];
        eta_sum[14][3]  = eta_sum_out_tmp[14][3];
        eta_sum[14][4]  = eta_sum_out_tmp[14][4];
        eta_sum[14][5]  = eta_sum_out_tmp[14][5];
        eta_sum[14][6]  = eta_sum_out_tmp[14][6];
        eta_sum[14][7]  = eta_sum_out_tmp[14][7];
        eta_sum[14][8]  = eta_sum_out_tmp[14][8];
        eta_sum[14][9]  = eta_sum_out_tmp[14][9];
        eta_sum[14][10]  = eta_sum_out_tmp[14][10];
        eta_sum[14][11]  = eta_sum_out_tmp[14][11];
        eta_sum[14][12]  = eta_sum_out_tmp[14][12];
        eta_sum[14][13]  = eta_sum_out_tmp[14][13];
        eta_sum[14][14]  = eta_sum_out_tmp[14][14];
        eta_sum[14][15]  = eta_sum_out_tmp[14][15];
        eta_sum[14][16]  = eta_sum_out_tmp[14][16];
        eta_sum[14][17]  = eta_sum_out_tmp[14][17];
        eta_sum[14][18]  = eta_sum_out_tmp[14][18];
        eta_sum[14][19]  = eta_sum_out_tmp[14][19];
        eta_sum[14][20]  = eta_sum_out_tmp[14][20];
        eta_sum[14][21]  = eta_sum_out_tmp[14][21];
        eta_sum[14][22]  = eta_sum_out_tmp[14][22];
        eta_sum[14][23]  = eta_sum_out_tmp[14][23];
        eta_sum[14][24]  = eta_sum_out_tmp[14][24];
        eta_sum[14][25]  = eta_sum_out_tmp[14][25];
        eta_sum[14][26]  = eta_sum_out_tmp[14][26];
        eta_sum[14][27]  = eta_sum_out_tmp[14][27];
        eta_sum[14][28]  = eta_sum_out_tmp[14][28];
        eta_sum[14][29]  = eta_sum_out_tmp[14][29];
        eta_sum[14][30]  = eta_sum_out_tmp[14][30];
        eta_sum[14][31]  = eta_sum_out_tmp[14][31];
        eta_sum[14][32]  = eta_sum_out_tmp[14][32];
        eta_sum[14][33]  = eta_sum_out_tmp[14][33];
        eta_sum[14][34]  = eta_sum_out_tmp[14][34];
        eta_sum[14][35]  = eta_sum_out_tmp[14][35];
        eta_sum[14][36]  = eta_sum_out_tmp[14][36];
        eta_sum[14][37]  = eta_sum_out_tmp[14][37];
        eta_sum[14][38]  = eta_sum_out_tmp[14][38];
        eta_sum[14][39]  = eta_sum_out_tmp[14][39];
        eta_sum[14][40]  = eta_sum_out_tmp[14][40];
        eta_sum[14][41]  = eta_sum_out_tmp[14][41];
    end
 
    6:begin 
        eta_sum[14][13]  = eta_sum_out_tmp[14][0];
        eta_sum[14][14]  = eta_sum_out_tmp[14][1];
        eta_sum[14][15]  = eta_sum_out_tmp[14][2];
        eta_sum[14][16]  = eta_sum_out_tmp[14][3];
        eta_sum[14][17]  = eta_sum_out_tmp[14][4];
        eta_sum[14][18]  = eta_sum_out_tmp[14][5];
        eta_sum[14][19]  = eta_sum_out_tmp[14][6];
        eta_sum[14][20]  = eta_sum_out_tmp[14][7];
        eta_sum[14][21]  = eta_sum_out_tmp[14][8];
        eta_sum[14][22]  = eta_sum_out_tmp[14][9];
        eta_sum[14][23]  = eta_sum_out_tmp[14][10];
        eta_sum[14][24]  = eta_sum_out_tmp[14][11];
        eta_sum[14][25]  = eta_sum_out_tmp[14][12];
        eta_sum[14][26]  = eta_sum_out_tmp[14][13];
        eta_sum[14][27]  = eta_sum_out_tmp[14][14];
        eta_sum[14][28]  = eta_sum_out_tmp[14][15];
        eta_sum[14][29]  = eta_sum_out_tmp[14][16];
        eta_sum[14][30]  = eta_sum_out_tmp[14][17];
        eta_sum[14][31]  = eta_sum_out_tmp[14][18];
        eta_sum[14][32]  = eta_sum_out_tmp[14][19];
        eta_sum[14][33]  = eta_sum_out_tmp[14][20];
        eta_sum[14][34]  = eta_sum_out_tmp[14][21];
        eta_sum[14][35]  = eta_sum_out_tmp[14][22];
        eta_sum[14][36]  = eta_sum_out_tmp[14][23];
        eta_sum[14][37]  = eta_sum_out_tmp[14][24];
        eta_sum[14][38]  = eta_sum_out_tmp[14][25];
        eta_sum[14][39]  = eta_sum_out_tmp[14][26];
        eta_sum[14][40]  = eta_sum_out_tmp[14][27];
        eta_sum[14][41]  = eta_sum_out_tmp[14][28];
        eta_sum[14][0]  = eta_sum_out_tmp[14][29];
        eta_sum[14][1]  = eta_sum_out_tmp[14][30];
        eta_sum[14][2]  = eta_sum_out_tmp[14][31];
        eta_sum[14][3]  = eta_sum_out_tmp[14][32];
        eta_sum[14][4]  = eta_sum_out_tmp[14][33];
        eta_sum[14][5]  = eta_sum_out_tmp[14][34];
        eta_sum[14][6]  = eta_sum_out_tmp[14][35];
        eta_sum[14][7]  = eta_sum_out_tmp[14][36];
        eta_sum[14][8]  = eta_sum_out_tmp[14][37];
        eta_sum[14][9]  = eta_sum_out_tmp[14][38];
        eta_sum[14][10]  = eta_sum_out_tmp[14][39];
        eta_sum[14][11]  = eta_sum_out_tmp[14][40];
        eta_sum[14][12]  = eta_sum_out_tmp[14][41];
    end
 
    7:begin 
        eta_sum[14][22]  = eta_sum_out_tmp[14][0];
        eta_sum[14][23]  = eta_sum_out_tmp[14][1];
        eta_sum[14][24]  = eta_sum_out_tmp[14][2];
        eta_sum[14][25]  = eta_sum_out_tmp[14][3];
        eta_sum[14][26]  = eta_sum_out_tmp[14][4];
        eta_sum[14][27]  = eta_sum_out_tmp[14][5];
        eta_sum[14][28]  = eta_sum_out_tmp[14][6];
        eta_sum[14][29]  = eta_sum_out_tmp[14][7];
        eta_sum[14][30]  = eta_sum_out_tmp[14][8];
        eta_sum[14][31]  = eta_sum_out_tmp[14][9];
        eta_sum[14][32]  = eta_sum_out_tmp[14][10];
        eta_sum[14][33]  = eta_sum_out_tmp[14][11];
        eta_sum[14][34]  = eta_sum_out_tmp[14][12];
        eta_sum[14][35]  = eta_sum_out_tmp[14][13];
        eta_sum[14][36]  = eta_sum_out_tmp[14][14];
        eta_sum[14][37]  = eta_sum_out_tmp[14][15];
        eta_sum[14][38]  = eta_sum_out_tmp[14][16];
        eta_sum[14][39]  = eta_sum_out_tmp[14][17];
        eta_sum[14][40]  = eta_sum_out_tmp[14][18];
        eta_sum[14][41]  = eta_sum_out_tmp[14][19];
        eta_sum[14][0]  = eta_sum_out_tmp[14][20];
        eta_sum[14][1]  = eta_sum_out_tmp[14][21];
        eta_sum[14][2]  = eta_sum_out_tmp[14][22];
        eta_sum[14][3]  = eta_sum_out_tmp[14][23];
        eta_sum[14][4]  = eta_sum_out_tmp[14][24];
        eta_sum[14][5]  = eta_sum_out_tmp[14][25];
        eta_sum[14][6]  = eta_sum_out_tmp[14][26];
        eta_sum[14][7]  = eta_sum_out_tmp[14][27];
        eta_sum[14][8]  = eta_sum_out_tmp[14][28];
        eta_sum[14][9]  = eta_sum_out_tmp[14][29];
        eta_sum[14][10]  = eta_sum_out_tmp[14][30];
        eta_sum[14][11]  = eta_sum_out_tmp[14][31];
        eta_sum[14][12]  = eta_sum_out_tmp[14][32];
        eta_sum[14][13]  = eta_sum_out_tmp[14][33];
        eta_sum[14][14]  = eta_sum_out_tmp[14][34];
        eta_sum[14][15]  = eta_sum_out_tmp[14][35];
        eta_sum[14][16]  = eta_sum_out_tmp[14][36];
        eta_sum[14][17]  = eta_sum_out_tmp[14][37];
        eta_sum[14][18]  = eta_sum_out_tmp[14][38];
        eta_sum[14][19]  = eta_sum_out_tmp[14][39];
        eta_sum[14][20]  = eta_sum_out_tmp[14][40];
        eta_sum[14][21]  = eta_sum_out_tmp[14][41];
    end
 
endcase
end

if (chk_n_output_valid[0] & active_cols[15]) begin
case (curr_layer)
    0:begin 
        eta_sum[15][0]  = eta_sum_out_tmp[15][0];
        eta_sum[15][1]  = eta_sum_out_tmp[15][1];
        eta_sum[15][2]  = eta_sum_out_tmp[15][2];
        eta_sum[15][3]  = eta_sum_out_tmp[15][3];
        eta_sum[15][4]  = eta_sum_out_tmp[15][4];
        eta_sum[15][5]  = eta_sum_out_tmp[15][5];
        eta_sum[15][6]  = eta_sum_out_tmp[15][6];
        eta_sum[15][7]  = eta_sum_out_tmp[15][7];
        eta_sum[15][8]  = eta_sum_out_tmp[15][8];
        eta_sum[15][9]  = eta_sum_out_tmp[15][9];
        eta_sum[15][10]  = eta_sum_out_tmp[15][10];
        eta_sum[15][11]  = eta_sum_out_tmp[15][11];
        eta_sum[15][12]  = eta_sum_out_tmp[15][12];
        eta_sum[15][13]  = eta_sum_out_tmp[15][13];
        eta_sum[15][14]  = eta_sum_out_tmp[15][14];
        eta_sum[15][15]  = eta_sum_out_tmp[15][15];
        eta_sum[15][16]  = eta_sum_out_tmp[15][16];
        eta_sum[15][17]  = eta_sum_out_tmp[15][17];
        eta_sum[15][18]  = eta_sum_out_tmp[15][18];
        eta_sum[15][19]  = eta_sum_out_tmp[15][19];
        eta_sum[15][20]  = eta_sum_out_tmp[15][20];
        eta_sum[15][21]  = eta_sum_out_tmp[15][21];
        eta_sum[15][22]  = eta_sum_out_tmp[15][22];
        eta_sum[15][23]  = eta_sum_out_tmp[15][23];
        eta_sum[15][24]  = eta_sum_out_tmp[15][24];
        eta_sum[15][25]  = eta_sum_out_tmp[15][25];
        eta_sum[15][26]  = eta_sum_out_tmp[15][26];
        eta_sum[15][27]  = eta_sum_out_tmp[15][27];
        eta_sum[15][28]  = eta_sum_out_tmp[15][28];
        eta_sum[15][29]  = eta_sum_out_tmp[15][29];
        eta_sum[15][30]  = eta_sum_out_tmp[15][30];
        eta_sum[15][31]  = eta_sum_out_tmp[15][31];
        eta_sum[15][32]  = eta_sum_out_tmp[15][32];
        eta_sum[15][33]  = eta_sum_out_tmp[15][33];
        eta_sum[15][34]  = eta_sum_out_tmp[15][34];
        eta_sum[15][35]  = eta_sum_out_tmp[15][35];
        eta_sum[15][36]  = eta_sum_out_tmp[15][36];
        eta_sum[15][37]  = eta_sum_out_tmp[15][37];
        eta_sum[15][38]  = eta_sum_out_tmp[15][38];
        eta_sum[15][39]  = eta_sum_out_tmp[15][39];
        eta_sum[15][40]  = eta_sum_out_tmp[15][40];
        eta_sum[15][41]  = eta_sum_out_tmp[15][41];
    end
 
    1:begin 
        eta_sum[15][0]  = eta_sum_out_tmp[15][0];
        eta_sum[15][1]  = eta_sum_out_tmp[15][1];
        eta_sum[15][2]  = eta_sum_out_tmp[15][2];
        eta_sum[15][3]  = eta_sum_out_tmp[15][3];
        eta_sum[15][4]  = eta_sum_out_tmp[15][4];
        eta_sum[15][5]  = eta_sum_out_tmp[15][5];
        eta_sum[15][6]  = eta_sum_out_tmp[15][6];
        eta_sum[15][7]  = eta_sum_out_tmp[15][7];
        eta_sum[15][8]  = eta_sum_out_tmp[15][8];
        eta_sum[15][9]  = eta_sum_out_tmp[15][9];
        eta_sum[15][10]  = eta_sum_out_tmp[15][10];
        eta_sum[15][11]  = eta_sum_out_tmp[15][11];
        eta_sum[15][12]  = eta_sum_out_tmp[15][12];
        eta_sum[15][13]  = eta_sum_out_tmp[15][13];
        eta_sum[15][14]  = eta_sum_out_tmp[15][14];
        eta_sum[15][15]  = eta_sum_out_tmp[15][15];
        eta_sum[15][16]  = eta_sum_out_tmp[15][16];
        eta_sum[15][17]  = eta_sum_out_tmp[15][17];
        eta_sum[15][18]  = eta_sum_out_tmp[15][18];
        eta_sum[15][19]  = eta_sum_out_tmp[15][19];
        eta_sum[15][20]  = eta_sum_out_tmp[15][20];
        eta_sum[15][21]  = eta_sum_out_tmp[15][21];
        eta_sum[15][22]  = eta_sum_out_tmp[15][22];
        eta_sum[15][23]  = eta_sum_out_tmp[15][23];
        eta_sum[15][24]  = eta_sum_out_tmp[15][24];
        eta_sum[15][25]  = eta_sum_out_tmp[15][25];
        eta_sum[15][26]  = eta_sum_out_tmp[15][26];
        eta_sum[15][27]  = eta_sum_out_tmp[15][27];
        eta_sum[15][28]  = eta_sum_out_tmp[15][28];
        eta_sum[15][29]  = eta_sum_out_tmp[15][29];
        eta_sum[15][30]  = eta_sum_out_tmp[15][30];
        eta_sum[15][31]  = eta_sum_out_tmp[15][31];
        eta_sum[15][32]  = eta_sum_out_tmp[15][32];
        eta_sum[15][33]  = eta_sum_out_tmp[15][33];
        eta_sum[15][34]  = eta_sum_out_tmp[15][34];
        eta_sum[15][35]  = eta_sum_out_tmp[15][35];
        eta_sum[15][36]  = eta_sum_out_tmp[15][36];
        eta_sum[15][37]  = eta_sum_out_tmp[15][37];
        eta_sum[15][38]  = eta_sum_out_tmp[15][38];
        eta_sum[15][39]  = eta_sum_out_tmp[15][39];
        eta_sum[15][40]  = eta_sum_out_tmp[15][40];
        eta_sum[15][41]  = eta_sum_out_tmp[15][41];
    end
 
    2:begin 
        eta_sum[15][0]  = eta_sum_out_tmp[15][0];
        eta_sum[15][1]  = eta_sum_out_tmp[15][1];
        eta_sum[15][2]  = eta_sum_out_tmp[15][2];
        eta_sum[15][3]  = eta_sum_out_tmp[15][3];
        eta_sum[15][4]  = eta_sum_out_tmp[15][4];
        eta_sum[15][5]  = eta_sum_out_tmp[15][5];
        eta_sum[15][6]  = eta_sum_out_tmp[15][6];
        eta_sum[15][7]  = eta_sum_out_tmp[15][7];
        eta_sum[15][8]  = eta_sum_out_tmp[15][8];
        eta_sum[15][9]  = eta_sum_out_tmp[15][9];
        eta_sum[15][10]  = eta_sum_out_tmp[15][10];
        eta_sum[15][11]  = eta_sum_out_tmp[15][11];
        eta_sum[15][12]  = eta_sum_out_tmp[15][12];
        eta_sum[15][13]  = eta_sum_out_tmp[15][13];
        eta_sum[15][14]  = eta_sum_out_tmp[15][14];
        eta_sum[15][15]  = eta_sum_out_tmp[15][15];
        eta_sum[15][16]  = eta_sum_out_tmp[15][16];
        eta_sum[15][17]  = eta_sum_out_tmp[15][17];
        eta_sum[15][18]  = eta_sum_out_tmp[15][18];
        eta_sum[15][19]  = eta_sum_out_tmp[15][19];
        eta_sum[15][20]  = eta_sum_out_tmp[15][20];
        eta_sum[15][21]  = eta_sum_out_tmp[15][21];
        eta_sum[15][22]  = eta_sum_out_tmp[15][22];
        eta_sum[15][23]  = eta_sum_out_tmp[15][23];
        eta_sum[15][24]  = eta_sum_out_tmp[15][24];
        eta_sum[15][25]  = eta_sum_out_tmp[15][25];
        eta_sum[15][26]  = eta_sum_out_tmp[15][26];
        eta_sum[15][27]  = eta_sum_out_tmp[15][27];
        eta_sum[15][28]  = eta_sum_out_tmp[15][28];
        eta_sum[15][29]  = eta_sum_out_tmp[15][29];
        eta_sum[15][30]  = eta_sum_out_tmp[15][30];
        eta_sum[15][31]  = eta_sum_out_tmp[15][31];
        eta_sum[15][32]  = eta_sum_out_tmp[15][32];
        eta_sum[15][33]  = eta_sum_out_tmp[15][33];
        eta_sum[15][34]  = eta_sum_out_tmp[15][34];
        eta_sum[15][35]  = eta_sum_out_tmp[15][35];
        eta_sum[15][36]  = eta_sum_out_tmp[15][36];
        eta_sum[15][37]  = eta_sum_out_tmp[15][37];
        eta_sum[15][38]  = eta_sum_out_tmp[15][38];
        eta_sum[15][39]  = eta_sum_out_tmp[15][39];
        eta_sum[15][40]  = eta_sum_out_tmp[15][40];
        eta_sum[15][41]  = eta_sum_out_tmp[15][41];
    end
 
    3:begin 
        eta_sum[15][0]  = eta_sum_out_tmp[15][0];
        eta_sum[15][1]  = eta_sum_out_tmp[15][1];
        eta_sum[15][2]  = eta_sum_out_tmp[15][2];
        eta_sum[15][3]  = eta_sum_out_tmp[15][3];
        eta_sum[15][4]  = eta_sum_out_tmp[15][4];
        eta_sum[15][5]  = eta_sum_out_tmp[15][5];
        eta_sum[15][6]  = eta_sum_out_tmp[15][6];
        eta_sum[15][7]  = eta_sum_out_tmp[15][7];
        eta_sum[15][8]  = eta_sum_out_tmp[15][8];
        eta_sum[15][9]  = eta_sum_out_tmp[15][9];
        eta_sum[15][10]  = eta_sum_out_tmp[15][10];
        eta_sum[15][11]  = eta_sum_out_tmp[15][11];
        eta_sum[15][12]  = eta_sum_out_tmp[15][12];
        eta_sum[15][13]  = eta_sum_out_tmp[15][13];
        eta_sum[15][14]  = eta_sum_out_tmp[15][14];
        eta_sum[15][15]  = eta_sum_out_tmp[15][15];
        eta_sum[15][16]  = eta_sum_out_tmp[15][16];
        eta_sum[15][17]  = eta_sum_out_tmp[15][17];
        eta_sum[15][18]  = eta_sum_out_tmp[15][18];
        eta_sum[15][19]  = eta_sum_out_tmp[15][19];
        eta_sum[15][20]  = eta_sum_out_tmp[15][20];
        eta_sum[15][21]  = eta_sum_out_tmp[15][21];
        eta_sum[15][22]  = eta_sum_out_tmp[15][22];
        eta_sum[15][23]  = eta_sum_out_tmp[15][23];
        eta_sum[15][24]  = eta_sum_out_tmp[15][24];
        eta_sum[15][25]  = eta_sum_out_tmp[15][25];
        eta_sum[15][26]  = eta_sum_out_tmp[15][26];
        eta_sum[15][27]  = eta_sum_out_tmp[15][27];
        eta_sum[15][28]  = eta_sum_out_tmp[15][28];
        eta_sum[15][29]  = eta_sum_out_tmp[15][29];
        eta_sum[15][30]  = eta_sum_out_tmp[15][30];
        eta_sum[15][31]  = eta_sum_out_tmp[15][31];
        eta_sum[15][32]  = eta_sum_out_tmp[15][32];
        eta_sum[15][33]  = eta_sum_out_tmp[15][33];
        eta_sum[15][34]  = eta_sum_out_tmp[15][34];
        eta_sum[15][35]  = eta_sum_out_tmp[15][35];
        eta_sum[15][36]  = eta_sum_out_tmp[15][36];
        eta_sum[15][37]  = eta_sum_out_tmp[15][37];
        eta_sum[15][38]  = eta_sum_out_tmp[15][38];
        eta_sum[15][39]  = eta_sum_out_tmp[15][39];
        eta_sum[15][40]  = eta_sum_out_tmp[15][40];
        eta_sum[15][41]  = eta_sum_out_tmp[15][41];
    end
 
    4:begin 
        eta_sum[15][0]  = eta_sum_out_tmp[15][0];
        eta_sum[15][1]  = eta_sum_out_tmp[15][1];
        eta_sum[15][2]  = eta_sum_out_tmp[15][2];
        eta_sum[15][3]  = eta_sum_out_tmp[15][3];
        eta_sum[15][4]  = eta_sum_out_tmp[15][4];
        eta_sum[15][5]  = eta_sum_out_tmp[15][5];
        eta_sum[15][6]  = eta_sum_out_tmp[15][6];
        eta_sum[15][7]  = eta_sum_out_tmp[15][7];
        eta_sum[15][8]  = eta_sum_out_tmp[15][8];
        eta_sum[15][9]  = eta_sum_out_tmp[15][9];
        eta_sum[15][10]  = eta_sum_out_tmp[15][10];
        eta_sum[15][11]  = eta_sum_out_tmp[15][11];
        eta_sum[15][12]  = eta_sum_out_tmp[15][12];
        eta_sum[15][13]  = eta_sum_out_tmp[15][13];
        eta_sum[15][14]  = eta_sum_out_tmp[15][14];
        eta_sum[15][15]  = eta_sum_out_tmp[15][15];
        eta_sum[15][16]  = eta_sum_out_tmp[15][16];
        eta_sum[15][17]  = eta_sum_out_tmp[15][17];
        eta_sum[15][18]  = eta_sum_out_tmp[15][18];
        eta_sum[15][19]  = eta_sum_out_tmp[15][19];
        eta_sum[15][20]  = eta_sum_out_tmp[15][20];
        eta_sum[15][21]  = eta_sum_out_tmp[15][21];
        eta_sum[15][22]  = eta_sum_out_tmp[15][22];
        eta_sum[15][23]  = eta_sum_out_tmp[15][23];
        eta_sum[15][24]  = eta_sum_out_tmp[15][24];
        eta_sum[15][25]  = eta_sum_out_tmp[15][25];
        eta_sum[15][26]  = eta_sum_out_tmp[15][26];
        eta_sum[15][27]  = eta_sum_out_tmp[15][27];
        eta_sum[15][28]  = eta_sum_out_tmp[15][28];
        eta_sum[15][29]  = eta_sum_out_tmp[15][29];
        eta_sum[15][30]  = eta_sum_out_tmp[15][30];
        eta_sum[15][31]  = eta_sum_out_tmp[15][31];
        eta_sum[15][32]  = eta_sum_out_tmp[15][32];
        eta_sum[15][33]  = eta_sum_out_tmp[15][33];
        eta_sum[15][34]  = eta_sum_out_tmp[15][34];
        eta_sum[15][35]  = eta_sum_out_tmp[15][35];
        eta_sum[15][36]  = eta_sum_out_tmp[15][36];
        eta_sum[15][37]  = eta_sum_out_tmp[15][37];
        eta_sum[15][38]  = eta_sum_out_tmp[15][38];
        eta_sum[15][39]  = eta_sum_out_tmp[15][39];
        eta_sum[15][40]  = eta_sum_out_tmp[15][40];
        eta_sum[15][41]  = eta_sum_out_tmp[15][41];
    end
 
    5:begin 
        eta_sum[15][0]  = eta_sum_out_tmp[15][0];
        eta_sum[15][1]  = eta_sum_out_tmp[15][1];
        eta_sum[15][2]  = eta_sum_out_tmp[15][2];
        eta_sum[15][3]  = eta_sum_out_tmp[15][3];
        eta_sum[15][4]  = eta_sum_out_tmp[15][4];
        eta_sum[15][5]  = eta_sum_out_tmp[15][5];
        eta_sum[15][6]  = eta_sum_out_tmp[15][6];
        eta_sum[15][7]  = eta_sum_out_tmp[15][7];
        eta_sum[15][8]  = eta_sum_out_tmp[15][8];
        eta_sum[15][9]  = eta_sum_out_tmp[15][9];
        eta_sum[15][10]  = eta_sum_out_tmp[15][10];
        eta_sum[15][11]  = eta_sum_out_tmp[15][11];
        eta_sum[15][12]  = eta_sum_out_tmp[15][12];
        eta_sum[15][13]  = eta_sum_out_tmp[15][13];
        eta_sum[15][14]  = eta_sum_out_tmp[15][14];
        eta_sum[15][15]  = eta_sum_out_tmp[15][15];
        eta_sum[15][16]  = eta_sum_out_tmp[15][16];
        eta_sum[15][17]  = eta_sum_out_tmp[15][17];
        eta_sum[15][18]  = eta_sum_out_tmp[15][18];
        eta_sum[15][19]  = eta_sum_out_tmp[15][19];
        eta_sum[15][20]  = eta_sum_out_tmp[15][20];
        eta_sum[15][21]  = eta_sum_out_tmp[15][21];
        eta_sum[15][22]  = eta_sum_out_tmp[15][22];
        eta_sum[15][23]  = eta_sum_out_tmp[15][23];
        eta_sum[15][24]  = eta_sum_out_tmp[15][24];
        eta_sum[15][25]  = eta_sum_out_tmp[15][25];
        eta_sum[15][26]  = eta_sum_out_tmp[15][26];
        eta_sum[15][27]  = eta_sum_out_tmp[15][27];
        eta_sum[15][28]  = eta_sum_out_tmp[15][28];
        eta_sum[15][29]  = eta_sum_out_tmp[15][29];
        eta_sum[15][30]  = eta_sum_out_tmp[15][30];
        eta_sum[15][31]  = eta_sum_out_tmp[15][31];
        eta_sum[15][32]  = eta_sum_out_tmp[15][32];
        eta_sum[15][33]  = eta_sum_out_tmp[15][33];
        eta_sum[15][34]  = eta_sum_out_tmp[15][34];
        eta_sum[15][35]  = eta_sum_out_tmp[15][35];
        eta_sum[15][36]  = eta_sum_out_tmp[15][36];
        eta_sum[15][37]  = eta_sum_out_tmp[15][37];
        eta_sum[15][38]  = eta_sum_out_tmp[15][38];
        eta_sum[15][39]  = eta_sum_out_tmp[15][39];
        eta_sum[15][40]  = eta_sum_out_tmp[15][40];
        eta_sum[15][41]  = eta_sum_out_tmp[15][41];
    end
 
    6:begin 
        eta_sum[15][0]  = eta_sum_out_tmp[15][0];
        eta_sum[15][1]  = eta_sum_out_tmp[15][1];
        eta_sum[15][2]  = eta_sum_out_tmp[15][2];
        eta_sum[15][3]  = eta_sum_out_tmp[15][3];
        eta_sum[15][4]  = eta_sum_out_tmp[15][4];
        eta_sum[15][5]  = eta_sum_out_tmp[15][5];
        eta_sum[15][6]  = eta_sum_out_tmp[15][6];
        eta_sum[15][7]  = eta_sum_out_tmp[15][7];
        eta_sum[15][8]  = eta_sum_out_tmp[15][8];
        eta_sum[15][9]  = eta_sum_out_tmp[15][9];
        eta_sum[15][10]  = eta_sum_out_tmp[15][10];
        eta_sum[15][11]  = eta_sum_out_tmp[15][11];
        eta_sum[15][12]  = eta_sum_out_tmp[15][12];
        eta_sum[15][13]  = eta_sum_out_tmp[15][13];
        eta_sum[15][14]  = eta_sum_out_tmp[15][14];
        eta_sum[15][15]  = eta_sum_out_tmp[15][15];
        eta_sum[15][16]  = eta_sum_out_tmp[15][16];
        eta_sum[15][17]  = eta_sum_out_tmp[15][17];
        eta_sum[15][18]  = eta_sum_out_tmp[15][18];
        eta_sum[15][19]  = eta_sum_out_tmp[15][19];
        eta_sum[15][20]  = eta_sum_out_tmp[15][20];
        eta_sum[15][21]  = eta_sum_out_tmp[15][21];
        eta_sum[15][22]  = eta_sum_out_tmp[15][22];
        eta_sum[15][23]  = eta_sum_out_tmp[15][23];
        eta_sum[15][24]  = eta_sum_out_tmp[15][24];
        eta_sum[15][25]  = eta_sum_out_tmp[15][25];
        eta_sum[15][26]  = eta_sum_out_tmp[15][26];
        eta_sum[15][27]  = eta_sum_out_tmp[15][27];
        eta_sum[15][28]  = eta_sum_out_tmp[15][28];
        eta_sum[15][29]  = eta_sum_out_tmp[15][29];
        eta_sum[15][30]  = eta_sum_out_tmp[15][30];
        eta_sum[15][31]  = eta_sum_out_tmp[15][31];
        eta_sum[15][32]  = eta_sum_out_tmp[15][32];
        eta_sum[15][33]  = eta_sum_out_tmp[15][33];
        eta_sum[15][34]  = eta_sum_out_tmp[15][34];
        eta_sum[15][35]  = eta_sum_out_tmp[15][35];
        eta_sum[15][36]  = eta_sum_out_tmp[15][36];
        eta_sum[15][37]  = eta_sum_out_tmp[15][37];
        eta_sum[15][38]  = eta_sum_out_tmp[15][38];
        eta_sum[15][39]  = eta_sum_out_tmp[15][39];
        eta_sum[15][40]  = eta_sum_out_tmp[15][40];
        eta_sum[15][41]  = eta_sum_out_tmp[15][41];
    end
 
    7:begin 
        eta_sum[15][24]  = eta_sum_out_tmp[15][0];
        eta_sum[15][25]  = eta_sum_out_tmp[15][1];
        eta_sum[15][26]  = eta_sum_out_tmp[15][2];
        eta_sum[15][27]  = eta_sum_out_tmp[15][3];
        eta_sum[15][28]  = eta_sum_out_tmp[15][4];
        eta_sum[15][29]  = eta_sum_out_tmp[15][5];
        eta_sum[15][30]  = eta_sum_out_tmp[15][6];
        eta_sum[15][31]  = eta_sum_out_tmp[15][7];
        eta_sum[15][32]  = eta_sum_out_tmp[15][8];
        eta_sum[15][33]  = eta_sum_out_tmp[15][9];
        eta_sum[15][34]  = eta_sum_out_tmp[15][10];
        eta_sum[15][35]  = eta_sum_out_tmp[15][11];
        eta_sum[15][36]  = eta_sum_out_tmp[15][12];
        eta_sum[15][37]  = eta_sum_out_tmp[15][13];
        eta_sum[15][38]  = eta_sum_out_tmp[15][14];
        eta_sum[15][39]  = eta_sum_out_tmp[15][15];
        eta_sum[15][40]  = eta_sum_out_tmp[15][16];
        eta_sum[15][41]  = eta_sum_out_tmp[15][17];
        eta_sum[15][0]  = eta_sum_out_tmp[15][18];
        eta_sum[15][1]  = eta_sum_out_tmp[15][19];
        eta_sum[15][2]  = eta_sum_out_tmp[15][20];
        eta_sum[15][3]  = eta_sum_out_tmp[15][21];
        eta_sum[15][4]  = eta_sum_out_tmp[15][22];
        eta_sum[15][5]  = eta_sum_out_tmp[15][23];
        eta_sum[15][6]  = eta_sum_out_tmp[15][24];
        eta_sum[15][7]  = eta_sum_out_tmp[15][25];
        eta_sum[15][8]  = eta_sum_out_tmp[15][26];
        eta_sum[15][9]  = eta_sum_out_tmp[15][27];
        eta_sum[15][10]  = eta_sum_out_tmp[15][28];
        eta_sum[15][11]  = eta_sum_out_tmp[15][29];
        eta_sum[15][12]  = eta_sum_out_tmp[15][30];
        eta_sum[15][13]  = eta_sum_out_tmp[15][31];
        eta_sum[15][14]  = eta_sum_out_tmp[15][32];
        eta_sum[15][15]  = eta_sum_out_tmp[15][33];
        eta_sum[15][16]  = eta_sum_out_tmp[15][34];
        eta_sum[15][17]  = eta_sum_out_tmp[15][35];
        eta_sum[15][18]  = eta_sum_out_tmp[15][36];
        eta_sum[15][19]  = eta_sum_out_tmp[15][37];
        eta_sum[15][20]  = eta_sum_out_tmp[15][38];
        eta_sum[15][21]  = eta_sum_out_tmp[15][39];
        eta_sum[15][22]  = eta_sum_out_tmp[15][40];
        eta_sum[15][23]  = eta_sum_out_tmp[15][41];
    end
 
endcase
end

end
