always @(posedge clk) begin 
if (chk_n_input_valid) begin
case (curr_layer)
    0:begin 
        llr_in_tmp[0][0]  = llr_new[0][40];
        llr_in_tmp[0][1]  = llr_new[0][41];
        llr_in_tmp[0][2]  = llr_new[0][0];
        llr_in_tmp[0][3]  = llr_new[0][1];
        llr_in_tmp[0][4]  = llr_new[0][2];
        llr_in_tmp[0][5]  = llr_new[0][3];
        llr_in_tmp[0][6]  = llr_new[0][4];
        llr_in_tmp[0][7]  = llr_new[0][5];
        llr_in_tmp[0][8]  = llr_new[0][6];
        llr_in_tmp[0][9]  = llr_new[0][7];
        llr_in_tmp[0][10]  = llr_new[0][8];
        llr_in_tmp[0][11]  = llr_new[0][9];
        llr_in_tmp[0][12]  = llr_new[0][10];
        llr_in_tmp[0][13]  = llr_new[0][11];
        llr_in_tmp[0][14]  = llr_new[0][12];
        llr_in_tmp[0][15]  = llr_new[0][13];
        llr_in_tmp[0][16]  = llr_new[0][14];
        llr_in_tmp[0][17]  = llr_new[0][15];
        llr_in_tmp[0][18]  = llr_new[0][16];
        llr_in_tmp[0][19]  = llr_new[0][17];
        llr_in_tmp[0][20]  = llr_new[0][18];
        llr_in_tmp[0][21]  = llr_new[0][19];
        llr_in_tmp[0][22]  = llr_new[0][20];
        llr_in_tmp[0][23]  = llr_new[0][21];
        llr_in_tmp[0][24]  = llr_new[0][22];
        llr_in_tmp[0][25]  = llr_new[0][23];
        llr_in_tmp[0][26]  = llr_new[0][24];
        llr_in_tmp[0][27]  = llr_new[0][25];
        llr_in_tmp[0][28]  = llr_new[0][26];
        llr_in_tmp[0][29]  = llr_new[0][27];
        llr_in_tmp[0][30]  = llr_new[0][28];
        llr_in_tmp[0][31]  = llr_new[0][29];
        llr_in_tmp[0][32]  = llr_new[0][30];
        llr_in_tmp[0][33]  = llr_new[0][31];
        llr_in_tmp[0][34]  = llr_new[0][32];
        llr_in_tmp[0][35]  = llr_new[0][33];
        llr_in_tmp[0][36]  = llr_new[0][34];
        llr_in_tmp[0][37]  = llr_new[0][35];
        llr_in_tmp[0][38]  = llr_new[0][36];
        llr_in_tmp[0][39]  = llr_new[0][37];
        llr_in_tmp[0][40]  = llr_new[0][38];
        llr_in_tmp[0][41]  = llr_new[0][39];
    end
 
    1:begin 
        llr_in_tmp[0][0]  = llr_new[0][34];
        llr_in_tmp[0][1]  = llr_new[0][35];
        llr_in_tmp[0][2]  = llr_new[0][36];
        llr_in_tmp[0][3]  = llr_new[0][37];
        llr_in_tmp[0][4]  = llr_new[0][38];
        llr_in_tmp[0][5]  = llr_new[0][39];
        llr_in_tmp[0][6]  = llr_new[0][40];
        llr_in_tmp[0][7]  = llr_new[0][41];
        llr_in_tmp[0][8]  = llr_new[0][0];
        llr_in_tmp[0][9]  = llr_new[0][1];
        llr_in_tmp[0][10]  = llr_new[0][2];
        llr_in_tmp[0][11]  = llr_new[0][3];
        llr_in_tmp[0][12]  = llr_new[0][4];
        llr_in_tmp[0][13]  = llr_new[0][5];
        llr_in_tmp[0][14]  = llr_new[0][6];
        llr_in_tmp[0][15]  = llr_new[0][7];
        llr_in_tmp[0][16]  = llr_new[0][8];
        llr_in_tmp[0][17]  = llr_new[0][9];
        llr_in_tmp[0][18]  = llr_new[0][10];
        llr_in_tmp[0][19]  = llr_new[0][11];
        llr_in_tmp[0][20]  = llr_new[0][12];
        llr_in_tmp[0][21]  = llr_new[0][13];
        llr_in_tmp[0][22]  = llr_new[0][14];
        llr_in_tmp[0][23]  = llr_new[0][15];
        llr_in_tmp[0][24]  = llr_new[0][16];
        llr_in_tmp[0][25]  = llr_new[0][17];
        llr_in_tmp[0][26]  = llr_new[0][18];
        llr_in_tmp[0][27]  = llr_new[0][19];
        llr_in_tmp[0][28]  = llr_new[0][20];
        llr_in_tmp[0][29]  = llr_new[0][21];
        llr_in_tmp[0][30]  = llr_new[0][22];
        llr_in_tmp[0][31]  = llr_new[0][23];
        llr_in_tmp[0][32]  = llr_new[0][24];
        llr_in_tmp[0][33]  = llr_new[0][25];
        llr_in_tmp[0][34]  = llr_new[0][26];
        llr_in_tmp[0][35]  = llr_new[0][27];
        llr_in_tmp[0][36]  = llr_new[0][28];
        llr_in_tmp[0][37]  = llr_new[0][29];
        llr_in_tmp[0][38]  = llr_new[0][30];
        llr_in_tmp[0][39]  = llr_new[0][31];
        llr_in_tmp[0][40]  = llr_new[0][32];
        llr_in_tmp[0][41]  = llr_new[0][33];
    end
 
    2:begin 
        llr_in_tmp[0][0]  = llr_new[0][0];
        llr_in_tmp[0][1]  = llr_new[0][1];
        llr_in_tmp[0][2]  = llr_new[0][2];
        llr_in_tmp[0][3]  = llr_new[0][3];
        llr_in_tmp[0][4]  = llr_new[0][4];
        llr_in_tmp[0][5]  = llr_new[0][5];
        llr_in_tmp[0][6]  = llr_new[0][6];
        llr_in_tmp[0][7]  = llr_new[0][7];
        llr_in_tmp[0][8]  = llr_new[0][8];
        llr_in_tmp[0][9]  = llr_new[0][9];
        llr_in_tmp[0][10]  = llr_new[0][10];
        llr_in_tmp[0][11]  = llr_new[0][11];
        llr_in_tmp[0][12]  = llr_new[0][12];
        llr_in_tmp[0][13]  = llr_new[0][13];
        llr_in_tmp[0][14]  = llr_new[0][14];
        llr_in_tmp[0][15]  = llr_new[0][15];
        llr_in_tmp[0][16]  = llr_new[0][16];
        llr_in_tmp[0][17]  = llr_new[0][17];
        llr_in_tmp[0][18]  = llr_new[0][18];
        llr_in_tmp[0][19]  = llr_new[0][19];
        llr_in_tmp[0][20]  = llr_new[0][20];
        llr_in_tmp[0][21]  = llr_new[0][21];
        llr_in_tmp[0][22]  = llr_new[0][22];
        llr_in_tmp[0][23]  = llr_new[0][23];
        llr_in_tmp[0][24]  = llr_new[0][24];
        llr_in_tmp[0][25]  = llr_new[0][25];
        llr_in_tmp[0][26]  = llr_new[0][26];
        llr_in_tmp[0][27]  = llr_new[0][27];
        llr_in_tmp[0][28]  = llr_new[0][28];
        llr_in_tmp[0][29]  = llr_new[0][29];
        llr_in_tmp[0][30]  = llr_new[0][30];
        llr_in_tmp[0][31]  = llr_new[0][31];
        llr_in_tmp[0][32]  = llr_new[0][32];
        llr_in_tmp[0][33]  = llr_new[0][33];
        llr_in_tmp[0][34]  = llr_new[0][34];
        llr_in_tmp[0][35]  = llr_new[0][35];
        llr_in_tmp[0][36]  = llr_new[0][36];
        llr_in_tmp[0][37]  = llr_new[0][37];
        llr_in_tmp[0][38]  = llr_new[0][38];
        llr_in_tmp[0][39]  = llr_new[0][39];
        llr_in_tmp[0][40]  = llr_new[0][40];
        llr_in_tmp[0][41]  = llr_new[0][41];
    end
 
    3:begin 
        llr_in_tmp[0][0]  = llr_new[0][0];
        llr_in_tmp[0][1]  = llr_new[0][1];
        llr_in_tmp[0][2]  = llr_new[0][2];
        llr_in_tmp[0][3]  = llr_new[0][3];
        llr_in_tmp[0][4]  = llr_new[0][4];
        llr_in_tmp[0][5]  = llr_new[0][5];
        llr_in_tmp[0][6]  = llr_new[0][6];
        llr_in_tmp[0][7]  = llr_new[0][7];
        llr_in_tmp[0][8]  = llr_new[0][8];
        llr_in_tmp[0][9]  = llr_new[0][9];
        llr_in_tmp[0][10]  = llr_new[0][10];
        llr_in_tmp[0][11]  = llr_new[0][11];
        llr_in_tmp[0][12]  = llr_new[0][12];
        llr_in_tmp[0][13]  = llr_new[0][13];
        llr_in_tmp[0][14]  = llr_new[0][14];
        llr_in_tmp[0][15]  = llr_new[0][15];
        llr_in_tmp[0][16]  = llr_new[0][16];
        llr_in_tmp[0][17]  = llr_new[0][17];
        llr_in_tmp[0][18]  = llr_new[0][18];
        llr_in_tmp[0][19]  = llr_new[0][19];
        llr_in_tmp[0][20]  = llr_new[0][20];
        llr_in_tmp[0][21]  = llr_new[0][21];
        llr_in_tmp[0][22]  = llr_new[0][22];
        llr_in_tmp[0][23]  = llr_new[0][23];
        llr_in_tmp[0][24]  = llr_new[0][24];
        llr_in_tmp[0][25]  = llr_new[0][25];
        llr_in_tmp[0][26]  = llr_new[0][26];
        llr_in_tmp[0][27]  = llr_new[0][27];
        llr_in_tmp[0][28]  = llr_new[0][28];
        llr_in_tmp[0][29]  = llr_new[0][29];
        llr_in_tmp[0][30]  = llr_new[0][30];
        llr_in_tmp[0][31]  = llr_new[0][31];
        llr_in_tmp[0][32]  = llr_new[0][32];
        llr_in_tmp[0][33]  = llr_new[0][33];
        llr_in_tmp[0][34]  = llr_new[0][34];
        llr_in_tmp[0][35]  = llr_new[0][35];
        llr_in_tmp[0][36]  = llr_new[0][36];
        llr_in_tmp[0][37]  = llr_new[0][37];
        llr_in_tmp[0][38]  = llr_new[0][38];
        llr_in_tmp[0][39]  = llr_new[0][39];
        llr_in_tmp[0][40]  = llr_new[0][40];
        llr_in_tmp[0][41]  = llr_new[0][41];
    end
 
    4:begin 
        llr_in_tmp[0][0]  = llr_new[0][35];
        llr_in_tmp[0][1]  = llr_new[0][36];
        llr_in_tmp[0][2]  = llr_new[0][37];
        llr_in_tmp[0][3]  = llr_new[0][38];
        llr_in_tmp[0][4]  = llr_new[0][39];
        llr_in_tmp[0][5]  = llr_new[0][40];
        llr_in_tmp[0][6]  = llr_new[0][41];
        llr_in_tmp[0][7]  = llr_new[0][0];
        llr_in_tmp[0][8]  = llr_new[0][1];
        llr_in_tmp[0][9]  = llr_new[0][2];
        llr_in_tmp[0][10]  = llr_new[0][3];
        llr_in_tmp[0][11]  = llr_new[0][4];
        llr_in_tmp[0][12]  = llr_new[0][5];
        llr_in_tmp[0][13]  = llr_new[0][6];
        llr_in_tmp[0][14]  = llr_new[0][7];
        llr_in_tmp[0][15]  = llr_new[0][8];
        llr_in_tmp[0][16]  = llr_new[0][9];
        llr_in_tmp[0][17]  = llr_new[0][10];
        llr_in_tmp[0][18]  = llr_new[0][11];
        llr_in_tmp[0][19]  = llr_new[0][12];
        llr_in_tmp[0][20]  = llr_new[0][13];
        llr_in_tmp[0][21]  = llr_new[0][14];
        llr_in_tmp[0][22]  = llr_new[0][15];
        llr_in_tmp[0][23]  = llr_new[0][16];
        llr_in_tmp[0][24]  = llr_new[0][17];
        llr_in_tmp[0][25]  = llr_new[0][18];
        llr_in_tmp[0][26]  = llr_new[0][19];
        llr_in_tmp[0][27]  = llr_new[0][20];
        llr_in_tmp[0][28]  = llr_new[0][21];
        llr_in_tmp[0][29]  = llr_new[0][22];
        llr_in_tmp[0][30]  = llr_new[0][23];
        llr_in_tmp[0][31]  = llr_new[0][24];
        llr_in_tmp[0][32]  = llr_new[0][25];
        llr_in_tmp[0][33]  = llr_new[0][26];
        llr_in_tmp[0][34]  = llr_new[0][27];
        llr_in_tmp[0][35]  = llr_new[0][28];
        llr_in_tmp[0][36]  = llr_new[0][29];
        llr_in_tmp[0][37]  = llr_new[0][30];
        llr_in_tmp[0][38]  = llr_new[0][31];
        llr_in_tmp[0][39]  = llr_new[0][32];
        llr_in_tmp[0][40]  = llr_new[0][33];
        llr_in_tmp[0][41]  = llr_new[0][34];
    end
 
    5:begin 
        llr_in_tmp[0][0]  = llr_new[0][29];
        llr_in_tmp[0][1]  = llr_new[0][30];
        llr_in_tmp[0][2]  = llr_new[0][31];
        llr_in_tmp[0][3]  = llr_new[0][32];
        llr_in_tmp[0][4]  = llr_new[0][33];
        llr_in_tmp[0][5]  = llr_new[0][34];
        llr_in_tmp[0][6]  = llr_new[0][35];
        llr_in_tmp[0][7]  = llr_new[0][36];
        llr_in_tmp[0][8]  = llr_new[0][37];
        llr_in_tmp[0][9]  = llr_new[0][38];
        llr_in_tmp[0][10]  = llr_new[0][39];
        llr_in_tmp[0][11]  = llr_new[0][40];
        llr_in_tmp[0][12]  = llr_new[0][41];
        llr_in_tmp[0][13]  = llr_new[0][0];
        llr_in_tmp[0][14]  = llr_new[0][1];
        llr_in_tmp[0][15]  = llr_new[0][2];
        llr_in_tmp[0][16]  = llr_new[0][3];
        llr_in_tmp[0][17]  = llr_new[0][4];
        llr_in_tmp[0][18]  = llr_new[0][5];
        llr_in_tmp[0][19]  = llr_new[0][6];
        llr_in_tmp[0][20]  = llr_new[0][7];
        llr_in_tmp[0][21]  = llr_new[0][8];
        llr_in_tmp[0][22]  = llr_new[0][9];
        llr_in_tmp[0][23]  = llr_new[0][10];
        llr_in_tmp[0][24]  = llr_new[0][11];
        llr_in_tmp[0][25]  = llr_new[0][12];
        llr_in_tmp[0][26]  = llr_new[0][13];
        llr_in_tmp[0][27]  = llr_new[0][14];
        llr_in_tmp[0][28]  = llr_new[0][15];
        llr_in_tmp[0][29]  = llr_new[0][16];
        llr_in_tmp[0][30]  = llr_new[0][17];
        llr_in_tmp[0][31]  = llr_new[0][18];
        llr_in_tmp[0][32]  = llr_new[0][19];
        llr_in_tmp[0][33]  = llr_new[0][20];
        llr_in_tmp[0][34]  = llr_new[0][21];
        llr_in_tmp[0][35]  = llr_new[0][22];
        llr_in_tmp[0][36]  = llr_new[0][23];
        llr_in_tmp[0][37]  = llr_new[0][24];
        llr_in_tmp[0][38]  = llr_new[0][25];
        llr_in_tmp[0][39]  = llr_new[0][26];
        llr_in_tmp[0][40]  = llr_new[0][27];
        llr_in_tmp[0][41]  = llr_new[0][28];
    end
 
    6:begin 
        llr_in_tmp[0][0]  = llr_new[0][0];
        llr_in_tmp[0][1]  = llr_new[0][1];
        llr_in_tmp[0][2]  = llr_new[0][2];
        llr_in_tmp[0][3]  = llr_new[0][3];
        llr_in_tmp[0][4]  = llr_new[0][4];
        llr_in_tmp[0][5]  = llr_new[0][5];
        llr_in_tmp[0][6]  = llr_new[0][6];
        llr_in_tmp[0][7]  = llr_new[0][7];
        llr_in_tmp[0][8]  = llr_new[0][8];
        llr_in_tmp[0][9]  = llr_new[0][9];
        llr_in_tmp[0][10]  = llr_new[0][10];
        llr_in_tmp[0][11]  = llr_new[0][11];
        llr_in_tmp[0][12]  = llr_new[0][12];
        llr_in_tmp[0][13]  = llr_new[0][13];
        llr_in_tmp[0][14]  = llr_new[0][14];
        llr_in_tmp[0][15]  = llr_new[0][15];
        llr_in_tmp[0][16]  = llr_new[0][16];
        llr_in_tmp[0][17]  = llr_new[0][17];
        llr_in_tmp[0][18]  = llr_new[0][18];
        llr_in_tmp[0][19]  = llr_new[0][19];
        llr_in_tmp[0][20]  = llr_new[0][20];
        llr_in_tmp[0][21]  = llr_new[0][21];
        llr_in_tmp[0][22]  = llr_new[0][22];
        llr_in_tmp[0][23]  = llr_new[0][23];
        llr_in_tmp[0][24]  = llr_new[0][24];
        llr_in_tmp[0][25]  = llr_new[0][25];
        llr_in_tmp[0][26]  = llr_new[0][26];
        llr_in_tmp[0][27]  = llr_new[0][27];
        llr_in_tmp[0][28]  = llr_new[0][28];
        llr_in_tmp[0][29]  = llr_new[0][29];
        llr_in_tmp[0][30]  = llr_new[0][30];
        llr_in_tmp[0][31]  = llr_new[0][31];
        llr_in_tmp[0][32]  = llr_new[0][32];
        llr_in_tmp[0][33]  = llr_new[0][33];
        llr_in_tmp[0][34]  = llr_new[0][34];
        llr_in_tmp[0][35]  = llr_new[0][35];
        llr_in_tmp[0][36]  = llr_new[0][36];
        llr_in_tmp[0][37]  = llr_new[0][37];
        llr_in_tmp[0][38]  = llr_new[0][38];
        llr_in_tmp[0][39]  = llr_new[0][39];
        llr_in_tmp[0][40]  = llr_new[0][40];
        llr_in_tmp[0][41]  = llr_new[0][41];
    end
 
    7:begin 
        llr_in_tmp[0][0]  = llr_new[0][0];
        llr_in_tmp[0][1]  = llr_new[0][1];
        llr_in_tmp[0][2]  = llr_new[0][2];
        llr_in_tmp[0][3]  = llr_new[0][3];
        llr_in_tmp[0][4]  = llr_new[0][4];
        llr_in_tmp[0][5]  = llr_new[0][5];
        llr_in_tmp[0][6]  = llr_new[0][6];
        llr_in_tmp[0][7]  = llr_new[0][7];
        llr_in_tmp[0][8]  = llr_new[0][8];
        llr_in_tmp[0][9]  = llr_new[0][9];
        llr_in_tmp[0][10]  = llr_new[0][10];
        llr_in_tmp[0][11]  = llr_new[0][11];
        llr_in_tmp[0][12]  = llr_new[0][12];
        llr_in_tmp[0][13]  = llr_new[0][13];
        llr_in_tmp[0][14]  = llr_new[0][14];
        llr_in_tmp[0][15]  = llr_new[0][15];
        llr_in_tmp[0][16]  = llr_new[0][16];
        llr_in_tmp[0][17]  = llr_new[0][17];
        llr_in_tmp[0][18]  = llr_new[0][18];
        llr_in_tmp[0][19]  = llr_new[0][19];
        llr_in_tmp[0][20]  = llr_new[0][20];
        llr_in_tmp[0][21]  = llr_new[0][21];
        llr_in_tmp[0][22]  = llr_new[0][22];
        llr_in_tmp[0][23]  = llr_new[0][23];
        llr_in_tmp[0][24]  = llr_new[0][24];
        llr_in_tmp[0][25]  = llr_new[0][25];
        llr_in_tmp[0][26]  = llr_new[0][26];
        llr_in_tmp[0][27]  = llr_new[0][27];
        llr_in_tmp[0][28]  = llr_new[0][28];
        llr_in_tmp[0][29]  = llr_new[0][29];
        llr_in_tmp[0][30]  = llr_new[0][30];
        llr_in_tmp[0][31]  = llr_new[0][31];
        llr_in_tmp[0][32]  = llr_new[0][32];
        llr_in_tmp[0][33]  = llr_new[0][33];
        llr_in_tmp[0][34]  = llr_new[0][34];
        llr_in_tmp[0][35]  = llr_new[0][35];
        llr_in_tmp[0][36]  = llr_new[0][36];
        llr_in_tmp[0][37]  = llr_new[0][37];
        llr_in_tmp[0][38]  = llr_new[0][38];
        llr_in_tmp[0][39]  = llr_new[0][39];
        llr_in_tmp[0][40]  = llr_new[0][40];
        llr_in_tmp[0][41]  = llr_new[0][41];
    end
 
endcase
end

if (chk_n_input_valid) begin
case (curr_layer)
    0:begin 
        llr_in_tmp[1][0]  = llr_new[1][0];
        llr_in_tmp[1][1]  = llr_new[1][1];
        llr_in_tmp[1][2]  = llr_new[1][2];
        llr_in_tmp[1][3]  = llr_new[1][3];
        llr_in_tmp[1][4]  = llr_new[1][4];
        llr_in_tmp[1][5]  = llr_new[1][5];
        llr_in_tmp[1][6]  = llr_new[1][6];
        llr_in_tmp[1][7]  = llr_new[1][7];
        llr_in_tmp[1][8]  = llr_new[1][8];
        llr_in_tmp[1][9]  = llr_new[1][9];
        llr_in_tmp[1][10]  = llr_new[1][10];
        llr_in_tmp[1][11]  = llr_new[1][11];
        llr_in_tmp[1][12]  = llr_new[1][12];
        llr_in_tmp[1][13]  = llr_new[1][13];
        llr_in_tmp[1][14]  = llr_new[1][14];
        llr_in_tmp[1][15]  = llr_new[1][15];
        llr_in_tmp[1][16]  = llr_new[1][16];
        llr_in_tmp[1][17]  = llr_new[1][17];
        llr_in_tmp[1][18]  = llr_new[1][18];
        llr_in_tmp[1][19]  = llr_new[1][19];
        llr_in_tmp[1][20]  = llr_new[1][20];
        llr_in_tmp[1][21]  = llr_new[1][21];
        llr_in_tmp[1][22]  = llr_new[1][22];
        llr_in_tmp[1][23]  = llr_new[1][23];
        llr_in_tmp[1][24]  = llr_new[1][24];
        llr_in_tmp[1][25]  = llr_new[1][25];
        llr_in_tmp[1][26]  = llr_new[1][26];
        llr_in_tmp[1][27]  = llr_new[1][27];
        llr_in_tmp[1][28]  = llr_new[1][28];
        llr_in_tmp[1][29]  = llr_new[1][29];
        llr_in_tmp[1][30]  = llr_new[1][30];
        llr_in_tmp[1][31]  = llr_new[1][31];
        llr_in_tmp[1][32]  = llr_new[1][32];
        llr_in_tmp[1][33]  = llr_new[1][33];
        llr_in_tmp[1][34]  = llr_new[1][34];
        llr_in_tmp[1][35]  = llr_new[1][35];
        llr_in_tmp[1][36]  = llr_new[1][36];
        llr_in_tmp[1][37]  = llr_new[1][37];
        llr_in_tmp[1][38]  = llr_new[1][38];
        llr_in_tmp[1][39]  = llr_new[1][39];
        llr_in_tmp[1][40]  = llr_new[1][40];
        llr_in_tmp[1][41]  = llr_new[1][41];
    end
 
    1:begin 
        llr_in_tmp[1][0]  = llr_new[1][0];
        llr_in_tmp[1][1]  = llr_new[1][1];
        llr_in_tmp[1][2]  = llr_new[1][2];
        llr_in_tmp[1][3]  = llr_new[1][3];
        llr_in_tmp[1][4]  = llr_new[1][4];
        llr_in_tmp[1][5]  = llr_new[1][5];
        llr_in_tmp[1][6]  = llr_new[1][6];
        llr_in_tmp[1][7]  = llr_new[1][7];
        llr_in_tmp[1][8]  = llr_new[1][8];
        llr_in_tmp[1][9]  = llr_new[1][9];
        llr_in_tmp[1][10]  = llr_new[1][10];
        llr_in_tmp[1][11]  = llr_new[1][11];
        llr_in_tmp[1][12]  = llr_new[1][12];
        llr_in_tmp[1][13]  = llr_new[1][13];
        llr_in_tmp[1][14]  = llr_new[1][14];
        llr_in_tmp[1][15]  = llr_new[1][15];
        llr_in_tmp[1][16]  = llr_new[1][16];
        llr_in_tmp[1][17]  = llr_new[1][17];
        llr_in_tmp[1][18]  = llr_new[1][18];
        llr_in_tmp[1][19]  = llr_new[1][19];
        llr_in_tmp[1][20]  = llr_new[1][20];
        llr_in_tmp[1][21]  = llr_new[1][21];
        llr_in_tmp[1][22]  = llr_new[1][22];
        llr_in_tmp[1][23]  = llr_new[1][23];
        llr_in_tmp[1][24]  = llr_new[1][24];
        llr_in_tmp[1][25]  = llr_new[1][25];
        llr_in_tmp[1][26]  = llr_new[1][26];
        llr_in_tmp[1][27]  = llr_new[1][27];
        llr_in_tmp[1][28]  = llr_new[1][28];
        llr_in_tmp[1][29]  = llr_new[1][29];
        llr_in_tmp[1][30]  = llr_new[1][30];
        llr_in_tmp[1][31]  = llr_new[1][31];
        llr_in_tmp[1][32]  = llr_new[1][32];
        llr_in_tmp[1][33]  = llr_new[1][33];
        llr_in_tmp[1][34]  = llr_new[1][34];
        llr_in_tmp[1][35]  = llr_new[1][35];
        llr_in_tmp[1][36]  = llr_new[1][36];
        llr_in_tmp[1][37]  = llr_new[1][37];
        llr_in_tmp[1][38]  = llr_new[1][38];
        llr_in_tmp[1][39]  = llr_new[1][39];
        llr_in_tmp[1][40]  = llr_new[1][40];
        llr_in_tmp[1][41]  = llr_new[1][41];
    end
 
    2:begin 
        llr_in_tmp[1][0]  = llr_new[1][36];
        llr_in_tmp[1][1]  = llr_new[1][37];
        llr_in_tmp[1][2]  = llr_new[1][38];
        llr_in_tmp[1][3]  = llr_new[1][39];
        llr_in_tmp[1][4]  = llr_new[1][40];
        llr_in_tmp[1][5]  = llr_new[1][41];
        llr_in_tmp[1][6]  = llr_new[1][0];
        llr_in_tmp[1][7]  = llr_new[1][1];
        llr_in_tmp[1][8]  = llr_new[1][2];
        llr_in_tmp[1][9]  = llr_new[1][3];
        llr_in_tmp[1][10]  = llr_new[1][4];
        llr_in_tmp[1][11]  = llr_new[1][5];
        llr_in_tmp[1][12]  = llr_new[1][6];
        llr_in_tmp[1][13]  = llr_new[1][7];
        llr_in_tmp[1][14]  = llr_new[1][8];
        llr_in_tmp[1][15]  = llr_new[1][9];
        llr_in_tmp[1][16]  = llr_new[1][10];
        llr_in_tmp[1][17]  = llr_new[1][11];
        llr_in_tmp[1][18]  = llr_new[1][12];
        llr_in_tmp[1][19]  = llr_new[1][13];
        llr_in_tmp[1][20]  = llr_new[1][14];
        llr_in_tmp[1][21]  = llr_new[1][15];
        llr_in_tmp[1][22]  = llr_new[1][16];
        llr_in_tmp[1][23]  = llr_new[1][17];
        llr_in_tmp[1][24]  = llr_new[1][18];
        llr_in_tmp[1][25]  = llr_new[1][19];
        llr_in_tmp[1][26]  = llr_new[1][20];
        llr_in_tmp[1][27]  = llr_new[1][21];
        llr_in_tmp[1][28]  = llr_new[1][22];
        llr_in_tmp[1][29]  = llr_new[1][23];
        llr_in_tmp[1][30]  = llr_new[1][24];
        llr_in_tmp[1][31]  = llr_new[1][25];
        llr_in_tmp[1][32]  = llr_new[1][26];
        llr_in_tmp[1][33]  = llr_new[1][27];
        llr_in_tmp[1][34]  = llr_new[1][28];
        llr_in_tmp[1][35]  = llr_new[1][29];
        llr_in_tmp[1][36]  = llr_new[1][30];
        llr_in_tmp[1][37]  = llr_new[1][31];
        llr_in_tmp[1][38]  = llr_new[1][32];
        llr_in_tmp[1][39]  = llr_new[1][33];
        llr_in_tmp[1][40]  = llr_new[1][34];
        llr_in_tmp[1][41]  = llr_new[1][35];
    end
 
    3:begin 
        llr_in_tmp[1][0]  = llr_new[1][27];
        llr_in_tmp[1][1]  = llr_new[1][28];
        llr_in_tmp[1][2]  = llr_new[1][29];
        llr_in_tmp[1][3]  = llr_new[1][30];
        llr_in_tmp[1][4]  = llr_new[1][31];
        llr_in_tmp[1][5]  = llr_new[1][32];
        llr_in_tmp[1][6]  = llr_new[1][33];
        llr_in_tmp[1][7]  = llr_new[1][34];
        llr_in_tmp[1][8]  = llr_new[1][35];
        llr_in_tmp[1][9]  = llr_new[1][36];
        llr_in_tmp[1][10]  = llr_new[1][37];
        llr_in_tmp[1][11]  = llr_new[1][38];
        llr_in_tmp[1][12]  = llr_new[1][39];
        llr_in_tmp[1][13]  = llr_new[1][40];
        llr_in_tmp[1][14]  = llr_new[1][41];
        llr_in_tmp[1][15]  = llr_new[1][0];
        llr_in_tmp[1][16]  = llr_new[1][1];
        llr_in_tmp[1][17]  = llr_new[1][2];
        llr_in_tmp[1][18]  = llr_new[1][3];
        llr_in_tmp[1][19]  = llr_new[1][4];
        llr_in_tmp[1][20]  = llr_new[1][5];
        llr_in_tmp[1][21]  = llr_new[1][6];
        llr_in_tmp[1][22]  = llr_new[1][7];
        llr_in_tmp[1][23]  = llr_new[1][8];
        llr_in_tmp[1][24]  = llr_new[1][9];
        llr_in_tmp[1][25]  = llr_new[1][10];
        llr_in_tmp[1][26]  = llr_new[1][11];
        llr_in_tmp[1][27]  = llr_new[1][12];
        llr_in_tmp[1][28]  = llr_new[1][13];
        llr_in_tmp[1][29]  = llr_new[1][14];
        llr_in_tmp[1][30]  = llr_new[1][15];
        llr_in_tmp[1][31]  = llr_new[1][16];
        llr_in_tmp[1][32]  = llr_new[1][17];
        llr_in_tmp[1][33]  = llr_new[1][18];
        llr_in_tmp[1][34]  = llr_new[1][19];
        llr_in_tmp[1][35]  = llr_new[1][20];
        llr_in_tmp[1][36]  = llr_new[1][21];
        llr_in_tmp[1][37]  = llr_new[1][22];
        llr_in_tmp[1][38]  = llr_new[1][23];
        llr_in_tmp[1][39]  = llr_new[1][24];
        llr_in_tmp[1][40]  = llr_new[1][25];
        llr_in_tmp[1][41]  = llr_new[1][26];
    end
 
    4:begin 
        llr_in_tmp[1][0]  = llr_new[1][0];
        llr_in_tmp[1][1]  = llr_new[1][1];
        llr_in_tmp[1][2]  = llr_new[1][2];
        llr_in_tmp[1][3]  = llr_new[1][3];
        llr_in_tmp[1][4]  = llr_new[1][4];
        llr_in_tmp[1][5]  = llr_new[1][5];
        llr_in_tmp[1][6]  = llr_new[1][6];
        llr_in_tmp[1][7]  = llr_new[1][7];
        llr_in_tmp[1][8]  = llr_new[1][8];
        llr_in_tmp[1][9]  = llr_new[1][9];
        llr_in_tmp[1][10]  = llr_new[1][10];
        llr_in_tmp[1][11]  = llr_new[1][11];
        llr_in_tmp[1][12]  = llr_new[1][12];
        llr_in_tmp[1][13]  = llr_new[1][13];
        llr_in_tmp[1][14]  = llr_new[1][14];
        llr_in_tmp[1][15]  = llr_new[1][15];
        llr_in_tmp[1][16]  = llr_new[1][16];
        llr_in_tmp[1][17]  = llr_new[1][17];
        llr_in_tmp[1][18]  = llr_new[1][18];
        llr_in_tmp[1][19]  = llr_new[1][19];
        llr_in_tmp[1][20]  = llr_new[1][20];
        llr_in_tmp[1][21]  = llr_new[1][21];
        llr_in_tmp[1][22]  = llr_new[1][22];
        llr_in_tmp[1][23]  = llr_new[1][23];
        llr_in_tmp[1][24]  = llr_new[1][24];
        llr_in_tmp[1][25]  = llr_new[1][25];
        llr_in_tmp[1][26]  = llr_new[1][26];
        llr_in_tmp[1][27]  = llr_new[1][27];
        llr_in_tmp[1][28]  = llr_new[1][28];
        llr_in_tmp[1][29]  = llr_new[1][29];
        llr_in_tmp[1][30]  = llr_new[1][30];
        llr_in_tmp[1][31]  = llr_new[1][31];
        llr_in_tmp[1][32]  = llr_new[1][32];
        llr_in_tmp[1][33]  = llr_new[1][33];
        llr_in_tmp[1][34]  = llr_new[1][34];
        llr_in_tmp[1][35]  = llr_new[1][35];
        llr_in_tmp[1][36]  = llr_new[1][36];
        llr_in_tmp[1][37]  = llr_new[1][37];
        llr_in_tmp[1][38]  = llr_new[1][38];
        llr_in_tmp[1][39]  = llr_new[1][39];
        llr_in_tmp[1][40]  = llr_new[1][40];
        llr_in_tmp[1][41]  = llr_new[1][41];
    end
 
    5:begin 
        llr_in_tmp[1][0]  = llr_new[1][0];
        llr_in_tmp[1][1]  = llr_new[1][1];
        llr_in_tmp[1][2]  = llr_new[1][2];
        llr_in_tmp[1][3]  = llr_new[1][3];
        llr_in_tmp[1][4]  = llr_new[1][4];
        llr_in_tmp[1][5]  = llr_new[1][5];
        llr_in_tmp[1][6]  = llr_new[1][6];
        llr_in_tmp[1][7]  = llr_new[1][7];
        llr_in_tmp[1][8]  = llr_new[1][8];
        llr_in_tmp[1][9]  = llr_new[1][9];
        llr_in_tmp[1][10]  = llr_new[1][10];
        llr_in_tmp[1][11]  = llr_new[1][11];
        llr_in_tmp[1][12]  = llr_new[1][12];
        llr_in_tmp[1][13]  = llr_new[1][13];
        llr_in_tmp[1][14]  = llr_new[1][14];
        llr_in_tmp[1][15]  = llr_new[1][15];
        llr_in_tmp[1][16]  = llr_new[1][16];
        llr_in_tmp[1][17]  = llr_new[1][17];
        llr_in_tmp[1][18]  = llr_new[1][18];
        llr_in_tmp[1][19]  = llr_new[1][19];
        llr_in_tmp[1][20]  = llr_new[1][20];
        llr_in_tmp[1][21]  = llr_new[1][21];
        llr_in_tmp[1][22]  = llr_new[1][22];
        llr_in_tmp[1][23]  = llr_new[1][23];
        llr_in_tmp[1][24]  = llr_new[1][24];
        llr_in_tmp[1][25]  = llr_new[1][25];
        llr_in_tmp[1][26]  = llr_new[1][26];
        llr_in_tmp[1][27]  = llr_new[1][27];
        llr_in_tmp[1][28]  = llr_new[1][28];
        llr_in_tmp[1][29]  = llr_new[1][29];
        llr_in_tmp[1][30]  = llr_new[1][30];
        llr_in_tmp[1][31]  = llr_new[1][31];
        llr_in_tmp[1][32]  = llr_new[1][32];
        llr_in_tmp[1][33]  = llr_new[1][33];
        llr_in_tmp[1][34]  = llr_new[1][34];
        llr_in_tmp[1][35]  = llr_new[1][35];
        llr_in_tmp[1][36]  = llr_new[1][36];
        llr_in_tmp[1][37]  = llr_new[1][37];
        llr_in_tmp[1][38]  = llr_new[1][38];
        llr_in_tmp[1][39]  = llr_new[1][39];
        llr_in_tmp[1][40]  = llr_new[1][40];
        llr_in_tmp[1][41]  = llr_new[1][41];
    end
 
    6:begin 
        llr_in_tmp[1][0]  = llr_new[1][31];
        llr_in_tmp[1][1]  = llr_new[1][32];
        llr_in_tmp[1][2]  = llr_new[1][33];
        llr_in_tmp[1][3]  = llr_new[1][34];
        llr_in_tmp[1][4]  = llr_new[1][35];
        llr_in_tmp[1][5]  = llr_new[1][36];
        llr_in_tmp[1][6]  = llr_new[1][37];
        llr_in_tmp[1][7]  = llr_new[1][38];
        llr_in_tmp[1][8]  = llr_new[1][39];
        llr_in_tmp[1][9]  = llr_new[1][40];
        llr_in_tmp[1][10]  = llr_new[1][41];
        llr_in_tmp[1][11]  = llr_new[1][0];
        llr_in_tmp[1][12]  = llr_new[1][1];
        llr_in_tmp[1][13]  = llr_new[1][2];
        llr_in_tmp[1][14]  = llr_new[1][3];
        llr_in_tmp[1][15]  = llr_new[1][4];
        llr_in_tmp[1][16]  = llr_new[1][5];
        llr_in_tmp[1][17]  = llr_new[1][6];
        llr_in_tmp[1][18]  = llr_new[1][7];
        llr_in_tmp[1][19]  = llr_new[1][8];
        llr_in_tmp[1][20]  = llr_new[1][9];
        llr_in_tmp[1][21]  = llr_new[1][10];
        llr_in_tmp[1][22]  = llr_new[1][11];
        llr_in_tmp[1][23]  = llr_new[1][12];
        llr_in_tmp[1][24]  = llr_new[1][13];
        llr_in_tmp[1][25]  = llr_new[1][14];
        llr_in_tmp[1][26]  = llr_new[1][15];
        llr_in_tmp[1][27]  = llr_new[1][16];
        llr_in_tmp[1][28]  = llr_new[1][17];
        llr_in_tmp[1][29]  = llr_new[1][18];
        llr_in_tmp[1][30]  = llr_new[1][19];
        llr_in_tmp[1][31]  = llr_new[1][20];
        llr_in_tmp[1][32]  = llr_new[1][21];
        llr_in_tmp[1][33]  = llr_new[1][22];
        llr_in_tmp[1][34]  = llr_new[1][23];
        llr_in_tmp[1][35]  = llr_new[1][24];
        llr_in_tmp[1][36]  = llr_new[1][25];
        llr_in_tmp[1][37]  = llr_new[1][26];
        llr_in_tmp[1][38]  = llr_new[1][27];
        llr_in_tmp[1][39]  = llr_new[1][28];
        llr_in_tmp[1][40]  = llr_new[1][29];
        llr_in_tmp[1][41]  = llr_new[1][30];
    end
 
    7:begin 
        llr_in_tmp[1][0]  = llr_new[1][22];
        llr_in_tmp[1][1]  = llr_new[1][23];
        llr_in_tmp[1][2]  = llr_new[1][24];
        llr_in_tmp[1][3]  = llr_new[1][25];
        llr_in_tmp[1][4]  = llr_new[1][26];
        llr_in_tmp[1][5]  = llr_new[1][27];
        llr_in_tmp[1][6]  = llr_new[1][28];
        llr_in_tmp[1][7]  = llr_new[1][29];
        llr_in_tmp[1][8]  = llr_new[1][30];
        llr_in_tmp[1][9]  = llr_new[1][31];
        llr_in_tmp[1][10]  = llr_new[1][32];
        llr_in_tmp[1][11]  = llr_new[1][33];
        llr_in_tmp[1][12]  = llr_new[1][34];
        llr_in_tmp[1][13]  = llr_new[1][35];
        llr_in_tmp[1][14]  = llr_new[1][36];
        llr_in_tmp[1][15]  = llr_new[1][37];
        llr_in_tmp[1][16]  = llr_new[1][38];
        llr_in_tmp[1][17]  = llr_new[1][39];
        llr_in_tmp[1][18]  = llr_new[1][40];
        llr_in_tmp[1][19]  = llr_new[1][41];
        llr_in_tmp[1][20]  = llr_new[1][0];
        llr_in_tmp[1][21]  = llr_new[1][1];
        llr_in_tmp[1][22]  = llr_new[1][2];
        llr_in_tmp[1][23]  = llr_new[1][3];
        llr_in_tmp[1][24]  = llr_new[1][4];
        llr_in_tmp[1][25]  = llr_new[1][5];
        llr_in_tmp[1][26]  = llr_new[1][6];
        llr_in_tmp[1][27]  = llr_new[1][7];
        llr_in_tmp[1][28]  = llr_new[1][8];
        llr_in_tmp[1][29]  = llr_new[1][9];
        llr_in_tmp[1][30]  = llr_new[1][10];
        llr_in_tmp[1][31]  = llr_new[1][11];
        llr_in_tmp[1][32]  = llr_new[1][12];
        llr_in_tmp[1][33]  = llr_new[1][13];
        llr_in_tmp[1][34]  = llr_new[1][14];
        llr_in_tmp[1][35]  = llr_new[1][15];
        llr_in_tmp[1][36]  = llr_new[1][16];
        llr_in_tmp[1][37]  = llr_new[1][17];
        llr_in_tmp[1][38]  = llr_new[1][18];
        llr_in_tmp[1][39]  = llr_new[1][19];
        llr_in_tmp[1][40]  = llr_new[1][20];
        llr_in_tmp[1][41]  = llr_new[1][21];
    end
 
endcase
end

if (chk_n_input_valid) begin
case (curr_layer)
    0:begin 
        llr_in_tmp[2][0]  = llr_new[2][38];
        llr_in_tmp[2][1]  = llr_new[2][39];
        llr_in_tmp[2][2]  = llr_new[2][40];
        llr_in_tmp[2][3]  = llr_new[2][41];
        llr_in_tmp[2][4]  = llr_new[2][0];
        llr_in_tmp[2][5]  = llr_new[2][1];
        llr_in_tmp[2][6]  = llr_new[2][2];
        llr_in_tmp[2][7]  = llr_new[2][3];
        llr_in_tmp[2][8]  = llr_new[2][4];
        llr_in_tmp[2][9]  = llr_new[2][5];
        llr_in_tmp[2][10]  = llr_new[2][6];
        llr_in_tmp[2][11]  = llr_new[2][7];
        llr_in_tmp[2][12]  = llr_new[2][8];
        llr_in_tmp[2][13]  = llr_new[2][9];
        llr_in_tmp[2][14]  = llr_new[2][10];
        llr_in_tmp[2][15]  = llr_new[2][11];
        llr_in_tmp[2][16]  = llr_new[2][12];
        llr_in_tmp[2][17]  = llr_new[2][13];
        llr_in_tmp[2][18]  = llr_new[2][14];
        llr_in_tmp[2][19]  = llr_new[2][15];
        llr_in_tmp[2][20]  = llr_new[2][16];
        llr_in_tmp[2][21]  = llr_new[2][17];
        llr_in_tmp[2][22]  = llr_new[2][18];
        llr_in_tmp[2][23]  = llr_new[2][19];
        llr_in_tmp[2][24]  = llr_new[2][20];
        llr_in_tmp[2][25]  = llr_new[2][21];
        llr_in_tmp[2][26]  = llr_new[2][22];
        llr_in_tmp[2][27]  = llr_new[2][23];
        llr_in_tmp[2][28]  = llr_new[2][24];
        llr_in_tmp[2][29]  = llr_new[2][25];
        llr_in_tmp[2][30]  = llr_new[2][26];
        llr_in_tmp[2][31]  = llr_new[2][27];
        llr_in_tmp[2][32]  = llr_new[2][28];
        llr_in_tmp[2][33]  = llr_new[2][29];
        llr_in_tmp[2][34]  = llr_new[2][30];
        llr_in_tmp[2][35]  = llr_new[2][31];
        llr_in_tmp[2][36]  = llr_new[2][32];
        llr_in_tmp[2][37]  = llr_new[2][33];
        llr_in_tmp[2][38]  = llr_new[2][34];
        llr_in_tmp[2][39]  = llr_new[2][35];
        llr_in_tmp[2][40]  = llr_new[2][36];
        llr_in_tmp[2][41]  = llr_new[2][37];
    end
 
    1:begin 
        llr_in_tmp[2][0]  = llr_new[2][35];
        llr_in_tmp[2][1]  = llr_new[2][36];
        llr_in_tmp[2][2]  = llr_new[2][37];
        llr_in_tmp[2][3]  = llr_new[2][38];
        llr_in_tmp[2][4]  = llr_new[2][39];
        llr_in_tmp[2][5]  = llr_new[2][40];
        llr_in_tmp[2][6]  = llr_new[2][41];
        llr_in_tmp[2][7]  = llr_new[2][0];
        llr_in_tmp[2][8]  = llr_new[2][1];
        llr_in_tmp[2][9]  = llr_new[2][2];
        llr_in_tmp[2][10]  = llr_new[2][3];
        llr_in_tmp[2][11]  = llr_new[2][4];
        llr_in_tmp[2][12]  = llr_new[2][5];
        llr_in_tmp[2][13]  = llr_new[2][6];
        llr_in_tmp[2][14]  = llr_new[2][7];
        llr_in_tmp[2][15]  = llr_new[2][8];
        llr_in_tmp[2][16]  = llr_new[2][9];
        llr_in_tmp[2][17]  = llr_new[2][10];
        llr_in_tmp[2][18]  = llr_new[2][11];
        llr_in_tmp[2][19]  = llr_new[2][12];
        llr_in_tmp[2][20]  = llr_new[2][13];
        llr_in_tmp[2][21]  = llr_new[2][14];
        llr_in_tmp[2][22]  = llr_new[2][15];
        llr_in_tmp[2][23]  = llr_new[2][16];
        llr_in_tmp[2][24]  = llr_new[2][17];
        llr_in_tmp[2][25]  = llr_new[2][18];
        llr_in_tmp[2][26]  = llr_new[2][19];
        llr_in_tmp[2][27]  = llr_new[2][20];
        llr_in_tmp[2][28]  = llr_new[2][21];
        llr_in_tmp[2][29]  = llr_new[2][22];
        llr_in_tmp[2][30]  = llr_new[2][23];
        llr_in_tmp[2][31]  = llr_new[2][24];
        llr_in_tmp[2][32]  = llr_new[2][25];
        llr_in_tmp[2][33]  = llr_new[2][26];
        llr_in_tmp[2][34]  = llr_new[2][27];
        llr_in_tmp[2][35]  = llr_new[2][28];
        llr_in_tmp[2][36]  = llr_new[2][29];
        llr_in_tmp[2][37]  = llr_new[2][30];
        llr_in_tmp[2][38]  = llr_new[2][31];
        llr_in_tmp[2][39]  = llr_new[2][32];
        llr_in_tmp[2][40]  = llr_new[2][33];
        llr_in_tmp[2][41]  = llr_new[2][34];
    end
 
    2:begin 
        llr_in_tmp[2][0]  = llr_new[2][0];
        llr_in_tmp[2][1]  = llr_new[2][1];
        llr_in_tmp[2][2]  = llr_new[2][2];
        llr_in_tmp[2][3]  = llr_new[2][3];
        llr_in_tmp[2][4]  = llr_new[2][4];
        llr_in_tmp[2][5]  = llr_new[2][5];
        llr_in_tmp[2][6]  = llr_new[2][6];
        llr_in_tmp[2][7]  = llr_new[2][7];
        llr_in_tmp[2][8]  = llr_new[2][8];
        llr_in_tmp[2][9]  = llr_new[2][9];
        llr_in_tmp[2][10]  = llr_new[2][10];
        llr_in_tmp[2][11]  = llr_new[2][11];
        llr_in_tmp[2][12]  = llr_new[2][12];
        llr_in_tmp[2][13]  = llr_new[2][13];
        llr_in_tmp[2][14]  = llr_new[2][14];
        llr_in_tmp[2][15]  = llr_new[2][15];
        llr_in_tmp[2][16]  = llr_new[2][16];
        llr_in_tmp[2][17]  = llr_new[2][17];
        llr_in_tmp[2][18]  = llr_new[2][18];
        llr_in_tmp[2][19]  = llr_new[2][19];
        llr_in_tmp[2][20]  = llr_new[2][20];
        llr_in_tmp[2][21]  = llr_new[2][21];
        llr_in_tmp[2][22]  = llr_new[2][22];
        llr_in_tmp[2][23]  = llr_new[2][23];
        llr_in_tmp[2][24]  = llr_new[2][24];
        llr_in_tmp[2][25]  = llr_new[2][25];
        llr_in_tmp[2][26]  = llr_new[2][26];
        llr_in_tmp[2][27]  = llr_new[2][27];
        llr_in_tmp[2][28]  = llr_new[2][28];
        llr_in_tmp[2][29]  = llr_new[2][29];
        llr_in_tmp[2][30]  = llr_new[2][30];
        llr_in_tmp[2][31]  = llr_new[2][31];
        llr_in_tmp[2][32]  = llr_new[2][32];
        llr_in_tmp[2][33]  = llr_new[2][33];
        llr_in_tmp[2][34]  = llr_new[2][34];
        llr_in_tmp[2][35]  = llr_new[2][35];
        llr_in_tmp[2][36]  = llr_new[2][36];
        llr_in_tmp[2][37]  = llr_new[2][37];
        llr_in_tmp[2][38]  = llr_new[2][38];
        llr_in_tmp[2][39]  = llr_new[2][39];
        llr_in_tmp[2][40]  = llr_new[2][40];
        llr_in_tmp[2][41]  = llr_new[2][41];
    end
 
    3:begin 
        llr_in_tmp[2][0]  = llr_new[2][0];
        llr_in_tmp[2][1]  = llr_new[2][1];
        llr_in_tmp[2][2]  = llr_new[2][2];
        llr_in_tmp[2][3]  = llr_new[2][3];
        llr_in_tmp[2][4]  = llr_new[2][4];
        llr_in_tmp[2][5]  = llr_new[2][5];
        llr_in_tmp[2][6]  = llr_new[2][6];
        llr_in_tmp[2][7]  = llr_new[2][7];
        llr_in_tmp[2][8]  = llr_new[2][8];
        llr_in_tmp[2][9]  = llr_new[2][9];
        llr_in_tmp[2][10]  = llr_new[2][10];
        llr_in_tmp[2][11]  = llr_new[2][11];
        llr_in_tmp[2][12]  = llr_new[2][12];
        llr_in_tmp[2][13]  = llr_new[2][13];
        llr_in_tmp[2][14]  = llr_new[2][14];
        llr_in_tmp[2][15]  = llr_new[2][15];
        llr_in_tmp[2][16]  = llr_new[2][16];
        llr_in_tmp[2][17]  = llr_new[2][17];
        llr_in_tmp[2][18]  = llr_new[2][18];
        llr_in_tmp[2][19]  = llr_new[2][19];
        llr_in_tmp[2][20]  = llr_new[2][20];
        llr_in_tmp[2][21]  = llr_new[2][21];
        llr_in_tmp[2][22]  = llr_new[2][22];
        llr_in_tmp[2][23]  = llr_new[2][23];
        llr_in_tmp[2][24]  = llr_new[2][24];
        llr_in_tmp[2][25]  = llr_new[2][25];
        llr_in_tmp[2][26]  = llr_new[2][26];
        llr_in_tmp[2][27]  = llr_new[2][27];
        llr_in_tmp[2][28]  = llr_new[2][28];
        llr_in_tmp[2][29]  = llr_new[2][29];
        llr_in_tmp[2][30]  = llr_new[2][30];
        llr_in_tmp[2][31]  = llr_new[2][31];
        llr_in_tmp[2][32]  = llr_new[2][32];
        llr_in_tmp[2][33]  = llr_new[2][33];
        llr_in_tmp[2][34]  = llr_new[2][34];
        llr_in_tmp[2][35]  = llr_new[2][35];
        llr_in_tmp[2][36]  = llr_new[2][36];
        llr_in_tmp[2][37]  = llr_new[2][37];
        llr_in_tmp[2][38]  = llr_new[2][38];
        llr_in_tmp[2][39]  = llr_new[2][39];
        llr_in_tmp[2][40]  = llr_new[2][40];
        llr_in_tmp[2][41]  = llr_new[2][41];
    end
 
    4:begin 
        llr_in_tmp[2][0]  = llr_new[2][41];
        llr_in_tmp[2][1]  = llr_new[2][0];
        llr_in_tmp[2][2]  = llr_new[2][1];
        llr_in_tmp[2][3]  = llr_new[2][2];
        llr_in_tmp[2][4]  = llr_new[2][3];
        llr_in_tmp[2][5]  = llr_new[2][4];
        llr_in_tmp[2][6]  = llr_new[2][5];
        llr_in_tmp[2][7]  = llr_new[2][6];
        llr_in_tmp[2][8]  = llr_new[2][7];
        llr_in_tmp[2][9]  = llr_new[2][8];
        llr_in_tmp[2][10]  = llr_new[2][9];
        llr_in_tmp[2][11]  = llr_new[2][10];
        llr_in_tmp[2][12]  = llr_new[2][11];
        llr_in_tmp[2][13]  = llr_new[2][12];
        llr_in_tmp[2][14]  = llr_new[2][13];
        llr_in_tmp[2][15]  = llr_new[2][14];
        llr_in_tmp[2][16]  = llr_new[2][15];
        llr_in_tmp[2][17]  = llr_new[2][16];
        llr_in_tmp[2][18]  = llr_new[2][17];
        llr_in_tmp[2][19]  = llr_new[2][18];
        llr_in_tmp[2][20]  = llr_new[2][19];
        llr_in_tmp[2][21]  = llr_new[2][20];
        llr_in_tmp[2][22]  = llr_new[2][21];
        llr_in_tmp[2][23]  = llr_new[2][22];
        llr_in_tmp[2][24]  = llr_new[2][23];
        llr_in_tmp[2][25]  = llr_new[2][24];
        llr_in_tmp[2][26]  = llr_new[2][25];
        llr_in_tmp[2][27]  = llr_new[2][26];
        llr_in_tmp[2][28]  = llr_new[2][27];
        llr_in_tmp[2][29]  = llr_new[2][28];
        llr_in_tmp[2][30]  = llr_new[2][29];
        llr_in_tmp[2][31]  = llr_new[2][30];
        llr_in_tmp[2][32]  = llr_new[2][31];
        llr_in_tmp[2][33]  = llr_new[2][32];
        llr_in_tmp[2][34]  = llr_new[2][33];
        llr_in_tmp[2][35]  = llr_new[2][34];
        llr_in_tmp[2][36]  = llr_new[2][35];
        llr_in_tmp[2][37]  = llr_new[2][36];
        llr_in_tmp[2][38]  = llr_new[2][37];
        llr_in_tmp[2][39]  = llr_new[2][38];
        llr_in_tmp[2][40]  = llr_new[2][39];
        llr_in_tmp[2][41]  = llr_new[2][40];
    end
 
    5:begin 
        llr_in_tmp[2][0]  = llr_new[2][0];
        llr_in_tmp[2][1]  = llr_new[2][1];
        llr_in_tmp[2][2]  = llr_new[2][2];
        llr_in_tmp[2][3]  = llr_new[2][3];
        llr_in_tmp[2][4]  = llr_new[2][4];
        llr_in_tmp[2][5]  = llr_new[2][5];
        llr_in_tmp[2][6]  = llr_new[2][6];
        llr_in_tmp[2][7]  = llr_new[2][7];
        llr_in_tmp[2][8]  = llr_new[2][8];
        llr_in_tmp[2][9]  = llr_new[2][9];
        llr_in_tmp[2][10]  = llr_new[2][10];
        llr_in_tmp[2][11]  = llr_new[2][11];
        llr_in_tmp[2][12]  = llr_new[2][12];
        llr_in_tmp[2][13]  = llr_new[2][13];
        llr_in_tmp[2][14]  = llr_new[2][14];
        llr_in_tmp[2][15]  = llr_new[2][15];
        llr_in_tmp[2][16]  = llr_new[2][16];
        llr_in_tmp[2][17]  = llr_new[2][17];
        llr_in_tmp[2][18]  = llr_new[2][18];
        llr_in_tmp[2][19]  = llr_new[2][19];
        llr_in_tmp[2][20]  = llr_new[2][20];
        llr_in_tmp[2][21]  = llr_new[2][21];
        llr_in_tmp[2][22]  = llr_new[2][22];
        llr_in_tmp[2][23]  = llr_new[2][23];
        llr_in_tmp[2][24]  = llr_new[2][24];
        llr_in_tmp[2][25]  = llr_new[2][25];
        llr_in_tmp[2][26]  = llr_new[2][26];
        llr_in_tmp[2][27]  = llr_new[2][27];
        llr_in_tmp[2][28]  = llr_new[2][28];
        llr_in_tmp[2][29]  = llr_new[2][29];
        llr_in_tmp[2][30]  = llr_new[2][30];
        llr_in_tmp[2][31]  = llr_new[2][31];
        llr_in_tmp[2][32]  = llr_new[2][32];
        llr_in_tmp[2][33]  = llr_new[2][33];
        llr_in_tmp[2][34]  = llr_new[2][34];
        llr_in_tmp[2][35]  = llr_new[2][35];
        llr_in_tmp[2][36]  = llr_new[2][36];
        llr_in_tmp[2][37]  = llr_new[2][37];
        llr_in_tmp[2][38]  = llr_new[2][38];
        llr_in_tmp[2][39]  = llr_new[2][39];
        llr_in_tmp[2][40]  = llr_new[2][40];
        llr_in_tmp[2][41]  = llr_new[2][41];
    end
 
    6:begin 
        llr_in_tmp[2][0]  = llr_new[2][0];
        llr_in_tmp[2][1]  = llr_new[2][1];
        llr_in_tmp[2][2]  = llr_new[2][2];
        llr_in_tmp[2][3]  = llr_new[2][3];
        llr_in_tmp[2][4]  = llr_new[2][4];
        llr_in_tmp[2][5]  = llr_new[2][5];
        llr_in_tmp[2][6]  = llr_new[2][6];
        llr_in_tmp[2][7]  = llr_new[2][7];
        llr_in_tmp[2][8]  = llr_new[2][8];
        llr_in_tmp[2][9]  = llr_new[2][9];
        llr_in_tmp[2][10]  = llr_new[2][10];
        llr_in_tmp[2][11]  = llr_new[2][11];
        llr_in_tmp[2][12]  = llr_new[2][12];
        llr_in_tmp[2][13]  = llr_new[2][13];
        llr_in_tmp[2][14]  = llr_new[2][14];
        llr_in_tmp[2][15]  = llr_new[2][15];
        llr_in_tmp[2][16]  = llr_new[2][16];
        llr_in_tmp[2][17]  = llr_new[2][17];
        llr_in_tmp[2][18]  = llr_new[2][18];
        llr_in_tmp[2][19]  = llr_new[2][19];
        llr_in_tmp[2][20]  = llr_new[2][20];
        llr_in_tmp[2][21]  = llr_new[2][21];
        llr_in_tmp[2][22]  = llr_new[2][22];
        llr_in_tmp[2][23]  = llr_new[2][23];
        llr_in_tmp[2][24]  = llr_new[2][24];
        llr_in_tmp[2][25]  = llr_new[2][25];
        llr_in_tmp[2][26]  = llr_new[2][26];
        llr_in_tmp[2][27]  = llr_new[2][27];
        llr_in_tmp[2][28]  = llr_new[2][28];
        llr_in_tmp[2][29]  = llr_new[2][29];
        llr_in_tmp[2][30]  = llr_new[2][30];
        llr_in_tmp[2][31]  = llr_new[2][31];
        llr_in_tmp[2][32]  = llr_new[2][32];
        llr_in_tmp[2][33]  = llr_new[2][33];
        llr_in_tmp[2][34]  = llr_new[2][34];
        llr_in_tmp[2][35]  = llr_new[2][35];
        llr_in_tmp[2][36]  = llr_new[2][36];
        llr_in_tmp[2][37]  = llr_new[2][37];
        llr_in_tmp[2][38]  = llr_new[2][38];
        llr_in_tmp[2][39]  = llr_new[2][39];
        llr_in_tmp[2][40]  = llr_new[2][40];
        llr_in_tmp[2][41]  = llr_new[2][41];
    end
 
    7:begin 
        llr_in_tmp[2][0]  = llr_new[2][0];
        llr_in_tmp[2][1]  = llr_new[2][1];
        llr_in_tmp[2][2]  = llr_new[2][2];
        llr_in_tmp[2][3]  = llr_new[2][3];
        llr_in_tmp[2][4]  = llr_new[2][4];
        llr_in_tmp[2][5]  = llr_new[2][5];
        llr_in_tmp[2][6]  = llr_new[2][6];
        llr_in_tmp[2][7]  = llr_new[2][7];
        llr_in_tmp[2][8]  = llr_new[2][8];
        llr_in_tmp[2][9]  = llr_new[2][9];
        llr_in_tmp[2][10]  = llr_new[2][10];
        llr_in_tmp[2][11]  = llr_new[2][11];
        llr_in_tmp[2][12]  = llr_new[2][12];
        llr_in_tmp[2][13]  = llr_new[2][13];
        llr_in_tmp[2][14]  = llr_new[2][14];
        llr_in_tmp[2][15]  = llr_new[2][15];
        llr_in_tmp[2][16]  = llr_new[2][16];
        llr_in_tmp[2][17]  = llr_new[2][17];
        llr_in_tmp[2][18]  = llr_new[2][18];
        llr_in_tmp[2][19]  = llr_new[2][19];
        llr_in_tmp[2][20]  = llr_new[2][20];
        llr_in_tmp[2][21]  = llr_new[2][21];
        llr_in_tmp[2][22]  = llr_new[2][22];
        llr_in_tmp[2][23]  = llr_new[2][23];
        llr_in_tmp[2][24]  = llr_new[2][24];
        llr_in_tmp[2][25]  = llr_new[2][25];
        llr_in_tmp[2][26]  = llr_new[2][26];
        llr_in_tmp[2][27]  = llr_new[2][27];
        llr_in_tmp[2][28]  = llr_new[2][28];
        llr_in_tmp[2][29]  = llr_new[2][29];
        llr_in_tmp[2][30]  = llr_new[2][30];
        llr_in_tmp[2][31]  = llr_new[2][31];
        llr_in_tmp[2][32]  = llr_new[2][32];
        llr_in_tmp[2][33]  = llr_new[2][33];
        llr_in_tmp[2][34]  = llr_new[2][34];
        llr_in_tmp[2][35]  = llr_new[2][35];
        llr_in_tmp[2][36]  = llr_new[2][36];
        llr_in_tmp[2][37]  = llr_new[2][37];
        llr_in_tmp[2][38]  = llr_new[2][38];
        llr_in_tmp[2][39]  = llr_new[2][39];
        llr_in_tmp[2][40]  = llr_new[2][40];
        llr_in_tmp[2][41]  = llr_new[2][41];
    end
 
endcase
end

if (chk_n_input_valid) begin
case (curr_layer)
    0:begin 
        llr_in_tmp[3][0]  = llr_new[3][0];
        llr_in_tmp[3][1]  = llr_new[3][1];
        llr_in_tmp[3][2]  = llr_new[3][2];
        llr_in_tmp[3][3]  = llr_new[3][3];
        llr_in_tmp[3][4]  = llr_new[3][4];
        llr_in_tmp[3][5]  = llr_new[3][5];
        llr_in_tmp[3][6]  = llr_new[3][6];
        llr_in_tmp[3][7]  = llr_new[3][7];
        llr_in_tmp[3][8]  = llr_new[3][8];
        llr_in_tmp[3][9]  = llr_new[3][9];
        llr_in_tmp[3][10]  = llr_new[3][10];
        llr_in_tmp[3][11]  = llr_new[3][11];
        llr_in_tmp[3][12]  = llr_new[3][12];
        llr_in_tmp[3][13]  = llr_new[3][13];
        llr_in_tmp[3][14]  = llr_new[3][14];
        llr_in_tmp[3][15]  = llr_new[3][15];
        llr_in_tmp[3][16]  = llr_new[3][16];
        llr_in_tmp[3][17]  = llr_new[3][17];
        llr_in_tmp[3][18]  = llr_new[3][18];
        llr_in_tmp[3][19]  = llr_new[3][19];
        llr_in_tmp[3][20]  = llr_new[3][20];
        llr_in_tmp[3][21]  = llr_new[3][21];
        llr_in_tmp[3][22]  = llr_new[3][22];
        llr_in_tmp[3][23]  = llr_new[3][23];
        llr_in_tmp[3][24]  = llr_new[3][24];
        llr_in_tmp[3][25]  = llr_new[3][25];
        llr_in_tmp[3][26]  = llr_new[3][26];
        llr_in_tmp[3][27]  = llr_new[3][27];
        llr_in_tmp[3][28]  = llr_new[3][28];
        llr_in_tmp[3][29]  = llr_new[3][29];
        llr_in_tmp[3][30]  = llr_new[3][30];
        llr_in_tmp[3][31]  = llr_new[3][31];
        llr_in_tmp[3][32]  = llr_new[3][32];
        llr_in_tmp[3][33]  = llr_new[3][33];
        llr_in_tmp[3][34]  = llr_new[3][34];
        llr_in_tmp[3][35]  = llr_new[3][35];
        llr_in_tmp[3][36]  = llr_new[3][36];
        llr_in_tmp[3][37]  = llr_new[3][37];
        llr_in_tmp[3][38]  = llr_new[3][38];
        llr_in_tmp[3][39]  = llr_new[3][39];
        llr_in_tmp[3][40]  = llr_new[3][40];
        llr_in_tmp[3][41]  = llr_new[3][41];
    end
 
    1:begin 
        llr_in_tmp[3][0]  = llr_new[3][0];
        llr_in_tmp[3][1]  = llr_new[3][1];
        llr_in_tmp[3][2]  = llr_new[3][2];
        llr_in_tmp[3][3]  = llr_new[3][3];
        llr_in_tmp[3][4]  = llr_new[3][4];
        llr_in_tmp[3][5]  = llr_new[3][5];
        llr_in_tmp[3][6]  = llr_new[3][6];
        llr_in_tmp[3][7]  = llr_new[3][7];
        llr_in_tmp[3][8]  = llr_new[3][8];
        llr_in_tmp[3][9]  = llr_new[3][9];
        llr_in_tmp[3][10]  = llr_new[3][10];
        llr_in_tmp[3][11]  = llr_new[3][11];
        llr_in_tmp[3][12]  = llr_new[3][12];
        llr_in_tmp[3][13]  = llr_new[3][13];
        llr_in_tmp[3][14]  = llr_new[3][14];
        llr_in_tmp[3][15]  = llr_new[3][15];
        llr_in_tmp[3][16]  = llr_new[3][16];
        llr_in_tmp[3][17]  = llr_new[3][17];
        llr_in_tmp[3][18]  = llr_new[3][18];
        llr_in_tmp[3][19]  = llr_new[3][19];
        llr_in_tmp[3][20]  = llr_new[3][20];
        llr_in_tmp[3][21]  = llr_new[3][21];
        llr_in_tmp[3][22]  = llr_new[3][22];
        llr_in_tmp[3][23]  = llr_new[3][23];
        llr_in_tmp[3][24]  = llr_new[3][24];
        llr_in_tmp[3][25]  = llr_new[3][25];
        llr_in_tmp[3][26]  = llr_new[3][26];
        llr_in_tmp[3][27]  = llr_new[3][27];
        llr_in_tmp[3][28]  = llr_new[3][28];
        llr_in_tmp[3][29]  = llr_new[3][29];
        llr_in_tmp[3][30]  = llr_new[3][30];
        llr_in_tmp[3][31]  = llr_new[3][31];
        llr_in_tmp[3][32]  = llr_new[3][32];
        llr_in_tmp[3][33]  = llr_new[3][33];
        llr_in_tmp[3][34]  = llr_new[3][34];
        llr_in_tmp[3][35]  = llr_new[3][35];
        llr_in_tmp[3][36]  = llr_new[3][36];
        llr_in_tmp[3][37]  = llr_new[3][37];
        llr_in_tmp[3][38]  = llr_new[3][38];
        llr_in_tmp[3][39]  = llr_new[3][39];
        llr_in_tmp[3][40]  = llr_new[3][40];
        llr_in_tmp[3][41]  = llr_new[3][41];
    end
 
    2:begin 
        llr_in_tmp[3][0]  = llr_new[3][31];
        llr_in_tmp[3][1]  = llr_new[3][32];
        llr_in_tmp[3][2]  = llr_new[3][33];
        llr_in_tmp[3][3]  = llr_new[3][34];
        llr_in_tmp[3][4]  = llr_new[3][35];
        llr_in_tmp[3][5]  = llr_new[3][36];
        llr_in_tmp[3][6]  = llr_new[3][37];
        llr_in_tmp[3][7]  = llr_new[3][38];
        llr_in_tmp[3][8]  = llr_new[3][39];
        llr_in_tmp[3][9]  = llr_new[3][40];
        llr_in_tmp[3][10]  = llr_new[3][41];
        llr_in_tmp[3][11]  = llr_new[3][0];
        llr_in_tmp[3][12]  = llr_new[3][1];
        llr_in_tmp[3][13]  = llr_new[3][2];
        llr_in_tmp[3][14]  = llr_new[3][3];
        llr_in_tmp[3][15]  = llr_new[3][4];
        llr_in_tmp[3][16]  = llr_new[3][5];
        llr_in_tmp[3][17]  = llr_new[3][6];
        llr_in_tmp[3][18]  = llr_new[3][7];
        llr_in_tmp[3][19]  = llr_new[3][8];
        llr_in_tmp[3][20]  = llr_new[3][9];
        llr_in_tmp[3][21]  = llr_new[3][10];
        llr_in_tmp[3][22]  = llr_new[3][11];
        llr_in_tmp[3][23]  = llr_new[3][12];
        llr_in_tmp[3][24]  = llr_new[3][13];
        llr_in_tmp[3][25]  = llr_new[3][14];
        llr_in_tmp[3][26]  = llr_new[3][15];
        llr_in_tmp[3][27]  = llr_new[3][16];
        llr_in_tmp[3][28]  = llr_new[3][17];
        llr_in_tmp[3][29]  = llr_new[3][18];
        llr_in_tmp[3][30]  = llr_new[3][19];
        llr_in_tmp[3][31]  = llr_new[3][20];
        llr_in_tmp[3][32]  = llr_new[3][21];
        llr_in_tmp[3][33]  = llr_new[3][22];
        llr_in_tmp[3][34]  = llr_new[3][23];
        llr_in_tmp[3][35]  = llr_new[3][24];
        llr_in_tmp[3][36]  = llr_new[3][25];
        llr_in_tmp[3][37]  = llr_new[3][26];
        llr_in_tmp[3][38]  = llr_new[3][27];
        llr_in_tmp[3][39]  = llr_new[3][28];
        llr_in_tmp[3][40]  = llr_new[3][29];
        llr_in_tmp[3][41]  = llr_new[3][30];
    end
 
    3:begin 
        llr_in_tmp[3][0]  = llr_new[3][18];
        llr_in_tmp[3][1]  = llr_new[3][19];
        llr_in_tmp[3][2]  = llr_new[3][20];
        llr_in_tmp[3][3]  = llr_new[3][21];
        llr_in_tmp[3][4]  = llr_new[3][22];
        llr_in_tmp[3][5]  = llr_new[3][23];
        llr_in_tmp[3][6]  = llr_new[3][24];
        llr_in_tmp[3][7]  = llr_new[3][25];
        llr_in_tmp[3][8]  = llr_new[3][26];
        llr_in_tmp[3][9]  = llr_new[3][27];
        llr_in_tmp[3][10]  = llr_new[3][28];
        llr_in_tmp[3][11]  = llr_new[3][29];
        llr_in_tmp[3][12]  = llr_new[3][30];
        llr_in_tmp[3][13]  = llr_new[3][31];
        llr_in_tmp[3][14]  = llr_new[3][32];
        llr_in_tmp[3][15]  = llr_new[3][33];
        llr_in_tmp[3][16]  = llr_new[3][34];
        llr_in_tmp[3][17]  = llr_new[3][35];
        llr_in_tmp[3][18]  = llr_new[3][36];
        llr_in_tmp[3][19]  = llr_new[3][37];
        llr_in_tmp[3][20]  = llr_new[3][38];
        llr_in_tmp[3][21]  = llr_new[3][39];
        llr_in_tmp[3][22]  = llr_new[3][40];
        llr_in_tmp[3][23]  = llr_new[3][41];
        llr_in_tmp[3][24]  = llr_new[3][0];
        llr_in_tmp[3][25]  = llr_new[3][1];
        llr_in_tmp[3][26]  = llr_new[3][2];
        llr_in_tmp[3][27]  = llr_new[3][3];
        llr_in_tmp[3][28]  = llr_new[3][4];
        llr_in_tmp[3][29]  = llr_new[3][5];
        llr_in_tmp[3][30]  = llr_new[3][6];
        llr_in_tmp[3][31]  = llr_new[3][7];
        llr_in_tmp[3][32]  = llr_new[3][8];
        llr_in_tmp[3][33]  = llr_new[3][9];
        llr_in_tmp[3][34]  = llr_new[3][10];
        llr_in_tmp[3][35]  = llr_new[3][11];
        llr_in_tmp[3][36]  = llr_new[3][12];
        llr_in_tmp[3][37]  = llr_new[3][13];
        llr_in_tmp[3][38]  = llr_new[3][14];
        llr_in_tmp[3][39]  = llr_new[3][15];
        llr_in_tmp[3][40]  = llr_new[3][16];
        llr_in_tmp[3][41]  = llr_new[3][17];
    end
 
    4:begin 
        llr_in_tmp[3][0]  = llr_new[3][0];
        llr_in_tmp[3][1]  = llr_new[3][1];
        llr_in_tmp[3][2]  = llr_new[3][2];
        llr_in_tmp[3][3]  = llr_new[3][3];
        llr_in_tmp[3][4]  = llr_new[3][4];
        llr_in_tmp[3][5]  = llr_new[3][5];
        llr_in_tmp[3][6]  = llr_new[3][6];
        llr_in_tmp[3][7]  = llr_new[3][7];
        llr_in_tmp[3][8]  = llr_new[3][8];
        llr_in_tmp[3][9]  = llr_new[3][9];
        llr_in_tmp[3][10]  = llr_new[3][10];
        llr_in_tmp[3][11]  = llr_new[3][11];
        llr_in_tmp[3][12]  = llr_new[3][12];
        llr_in_tmp[3][13]  = llr_new[3][13];
        llr_in_tmp[3][14]  = llr_new[3][14];
        llr_in_tmp[3][15]  = llr_new[3][15];
        llr_in_tmp[3][16]  = llr_new[3][16];
        llr_in_tmp[3][17]  = llr_new[3][17];
        llr_in_tmp[3][18]  = llr_new[3][18];
        llr_in_tmp[3][19]  = llr_new[3][19];
        llr_in_tmp[3][20]  = llr_new[3][20];
        llr_in_tmp[3][21]  = llr_new[3][21];
        llr_in_tmp[3][22]  = llr_new[3][22];
        llr_in_tmp[3][23]  = llr_new[3][23];
        llr_in_tmp[3][24]  = llr_new[3][24];
        llr_in_tmp[3][25]  = llr_new[3][25];
        llr_in_tmp[3][26]  = llr_new[3][26];
        llr_in_tmp[3][27]  = llr_new[3][27];
        llr_in_tmp[3][28]  = llr_new[3][28];
        llr_in_tmp[3][29]  = llr_new[3][29];
        llr_in_tmp[3][30]  = llr_new[3][30];
        llr_in_tmp[3][31]  = llr_new[3][31];
        llr_in_tmp[3][32]  = llr_new[3][32];
        llr_in_tmp[3][33]  = llr_new[3][33];
        llr_in_tmp[3][34]  = llr_new[3][34];
        llr_in_tmp[3][35]  = llr_new[3][35];
        llr_in_tmp[3][36]  = llr_new[3][36];
        llr_in_tmp[3][37]  = llr_new[3][37];
        llr_in_tmp[3][38]  = llr_new[3][38];
        llr_in_tmp[3][39]  = llr_new[3][39];
        llr_in_tmp[3][40]  = llr_new[3][40];
        llr_in_tmp[3][41]  = llr_new[3][41];
    end
 
    5:begin 
        llr_in_tmp[3][0]  = llr_new[3][0];
        llr_in_tmp[3][1]  = llr_new[3][1];
        llr_in_tmp[3][2]  = llr_new[3][2];
        llr_in_tmp[3][3]  = llr_new[3][3];
        llr_in_tmp[3][4]  = llr_new[3][4];
        llr_in_tmp[3][5]  = llr_new[3][5];
        llr_in_tmp[3][6]  = llr_new[3][6];
        llr_in_tmp[3][7]  = llr_new[3][7];
        llr_in_tmp[3][8]  = llr_new[3][8];
        llr_in_tmp[3][9]  = llr_new[3][9];
        llr_in_tmp[3][10]  = llr_new[3][10];
        llr_in_tmp[3][11]  = llr_new[3][11];
        llr_in_tmp[3][12]  = llr_new[3][12];
        llr_in_tmp[3][13]  = llr_new[3][13];
        llr_in_tmp[3][14]  = llr_new[3][14];
        llr_in_tmp[3][15]  = llr_new[3][15];
        llr_in_tmp[3][16]  = llr_new[3][16];
        llr_in_tmp[3][17]  = llr_new[3][17];
        llr_in_tmp[3][18]  = llr_new[3][18];
        llr_in_tmp[3][19]  = llr_new[3][19];
        llr_in_tmp[3][20]  = llr_new[3][20];
        llr_in_tmp[3][21]  = llr_new[3][21];
        llr_in_tmp[3][22]  = llr_new[3][22];
        llr_in_tmp[3][23]  = llr_new[3][23];
        llr_in_tmp[3][24]  = llr_new[3][24];
        llr_in_tmp[3][25]  = llr_new[3][25];
        llr_in_tmp[3][26]  = llr_new[3][26];
        llr_in_tmp[3][27]  = llr_new[3][27];
        llr_in_tmp[3][28]  = llr_new[3][28];
        llr_in_tmp[3][29]  = llr_new[3][29];
        llr_in_tmp[3][30]  = llr_new[3][30];
        llr_in_tmp[3][31]  = llr_new[3][31];
        llr_in_tmp[3][32]  = llr_new[3][32];
        llr_in_tmp[3][33]  = llr_new[3][33];
        llr_in_tmp[3][34]  = llr_new[3][34];
        llr_in_tmp[3][35]  = llr_new[3][35];
        llr_in_tmp[3][36]  = llr_new[3][36];
        llr_in_tmp[3][37]  = llr_new[3][37];
        llr_in_tmp[3][38]  = llr_new[3][38];
        llr_in_tmp[3][39]  = llr_new[3][39];
        llr_in_tmp[3][40]  = llr_new[3][40];
        llr_in_tmp[3][41]  = llr_new[3][41];
    end
 
    6:begin 
        llr_in_tmp[3][0]  = llr_new[3][23];
        llr_in_tmp[3][1]  = llr_new[3][24];
        llr_in_tmp[3][2]  = llr_new[3][25];
        llr_in_tmp[3][3]  = llr_new[3][26];
        llr_in_tmp[3][4]  = llr_new[3][27];
        llr_in_tmp[3][5]  = llr_new[3][28];
        llr_in_tmp[3][6]  = llr_new[3][29];
        llr_in_tmp[3][7]  = llr_new[3][30];
        llr_in_tmp[3][8]  = llr_new[3][31];
        llr_in_tmp[3][9]  = llr_new[3][32];
        llr_in_tmp[3][10]  = llr_new[3][33];
        llr_in_tmp[3][11]  = llr_new[3][34];
        llr_in_tmp[3][12]  = llr_new[3][35];
        llr_in_tmp[3][13]  = llr_new[3][36];
        llr_in_tmp[3][14]  = llr_new[3][37];
        llr_in_tmp[3][15]  = llr_new[3][38];
        llr_in_tmp[3][16]  = llr_new[3][39];
        llr_in_tmp[3][17]  = llr_new[3][40];
        llr_in_tmp[3][18]  = llr_new[3][41];
        llr_in_tmp[3][19]  = llr_new[3][0];
        llr_in_tmp[3][20]  = llr_new[3][1];
        llr_in_tmp[3][21]  = llr_new[3][2];
        llr_in_tmp[3][22]  = llr_new[3][3];
        llr_in_tmp[3][23]  = llr_new[3][4];
        llr_in_tmp[3][24]  = llr_new[3][5];
        llr_in_tmp[3][25]  = llr_new[3][6];
        llr_in_tmp[3][26]  = llr_new[3][7];
        llr_in_tmp[3][27]  = llr_new[3][8];
        llr_in_tmp[3][28]  = llr_new[3][9];
        llr_in_tmp[3][29]  = llr_new[3][10];
        llr_in_tmp[3][30]  = llr_new[3][11];
        llr_in_tmp[3][31]  = llr_new[3][12];
        llr_in_tmp[3][32]  = llr_new[3][13];
        llr_in_tmp[3][33]  = llr_new[3][14];
        llr_in_tmp[3][34]  = llr_new[3][15];
        llr_in_tmp[3][35]  = llr_new[3][16];
        llr_in_tmp[3][36]  = llr_new[3][17];
        llr_in_tmp[3][37]  = llr_new[3][18];
        llr_in_tmp[3][38]  = llr_new[3][19];
        llr_in_tmp[3][39]  = llr_new[3][20];
        llr_in_tmp[3][40]  = llr_new[3][21];
        llr_in_tmp[3][41]  = llr_new[3][22];
    end
 
    7:begin 
        llr_in_tmp[3][0]  = llr_new[3][34];
        llr_in_tmp[3][1]  = llr_new[3][35];
        llr_in_tmp[3][2]  = llr_new[3][36];
        llr_in_tmp[3][3]  = llr_new[3][37];
        llr_in_tmp[3][4]  = llr_new[3][38];
        llr_in_tmp[3][5]  = llr_new[3][39];
        llr_in_tmp[3][6]  = llr_new[3][40];
        llr_in_tmp[3][7]  = llr_new[3][41];
        llr_in_tmp[3][8]  = llr_new[3][0];
        llr_in_tmp[3][9]  = llr_new[3][1];
        llr_in_tmp[3][10]  = llr_new[3][2];
        llr_in_tmp[3][11]  = llr_new[3][3];
        llr_in_tmp[3][12]  = llr_new[3][4];
        llr_in_tmp[3][13]  = llr_new[3][5];
        llr_in_tmp[3][14]  = llr_new[3][6];
        llr_in_tmp[3][15]  = llr_new[3][7];
        llr_in_tmp[3][16]  = llr_new[3][8];
        llr_in_tmp[3][17]  = llr_new[3][9];
        llr_in_tmp[3][18]  = llr_new[3][10];
        llr_in_tmp[3][19]  = llr_new[3][11];
        llr_in_tmp[3][20]  = llr_new[3][12];
        llr_in_tmp[3][21]  = llr_new[3][13];
        llr_in_tmp[3][22]  = llr_new[3][14];
        llr_in_tmp[3][23]  = llr_new[3][15];
        llr_in_tmp[3][24]  = llr_new[3][16];
        llr_in_tmp[3][25]  = llr_new[3][17];
        llr_in_tmp[3][26]  = llr_new[3][18];
        llr_in_tmp[3][27]  = llr_new[3][19];
        llr_in_tmp[3][28]  = llr_new[3][20];
        llr_in_tmp[3][29]  = llr_new[3][21];
        llr_in_tmp[3][30]  = llr_new[3][22];
        llr_in_tmp[3][31]  = llr_new[3][23];
        llr_in_tmp[3][32]  = llr_new[3][24];
        llr_in_tmp[3][33]  = llr_new[3][25];
        llr_in_tmp[3][34]  = llr_new[3][26];
        llr_in_tmp[3][35]  = llr_new[3][27];
        llr_in_tmp[3][36]  = llr_new[3][28];
        llr_in_tmp[3][37]  = llr_new[3][29];
        llr_in_tmp[3][38]  = llr_new[3][30];
        llr_in_tmp[3][39]  = llr_new[3][31];
        llr_in_tmp[3][40]  = llr_new[3][32];
        llr_in_tmp[3][41]  = llr_new[3][33];
    end
 
endcase
end

if (chk_n_input_valid) begin
case (curr_layer)
    0:begin 
        llr_in_tmp[4][0]  = llr_new[4][13];
        llr_in_tmp[4][1]  = llr_new[4][14];
        llr_in_tmp[4][2]  = llr_new[4][15];
        llr_in_tmp[4][3]  = llr_new[4][16];
        llr_in_tmp[4][4]  = llr_new[4][17];
        llr_in_tmp[4][5]  = llr_new[4][18];
        llr_in_tmp[4][6]  = llr_new[4][19];
        llr_in_tmp[4][7]  = llr_new[4][20];
        llr_in_tmp[4][8]  = llr_new[4][21];
        llr_in_tmp[4][9]  = llr_new[4][22];
        llr_in_tmp[4][10]  = llr_new[4][23];
        llr_in_tmp[4][11]  = llr_new[4][24];
        llr_in_tmp[4][12]  = llr_new[4][25];
        llr_in_tmp[4][13]  = llr_new[4][26];
        llr_in_tmp[4][14]  = llr_new[4][27];
        llr_in_tmp[4][15]  = llr_new[4][28];
        llr_in_tmp[4][16]  = llr_new[4][29];
        llr_in_tmp[4][17]  = llr_new[4][30];
        llr_in_tmp[4][18]  = llr_new[4][31];
        llr_in_tmp[4][19]  = llr_new[4][32];
        llr_in_tmp[4][20]  = llr_new[4][33];
        llr_in_tmp[4][21]  = llr_new[4][34];
        llr_in_tmp[4][22]  = llr_new[4][35];
        llr_in_tmp[4][23]  = llr_new[4][36];
        llr_in_tmp[4][24]  = llr_new[4][37];
        llr_in_tmp[4][25]  = llr_new[4][38];
        llr_in_tmp[4][26]  = llr_new[4][39];
        llr_in_tmp[4][27]  = llr_new[4][40];
        llr_in_tmp[4][28]  = llr_new[4][41];
        llr_in_tmp[4][29]  = llr_new[4][0];
        llr_in_tmp[4][30]  = llr_new[4][1];
        llr_in_tmp[4][31]  = llr_new[4][2];
        llr_in_tmp[4][32]  = llr_new[4][3];
        llr_in_tmp[4][33]  = llr_new[4][4];
        llr_in_tmp[4][34]  = llr_new[4][5];
        llr_in_tmp[4][35]  = llr_new[4][6];
        llr_in_tmp[4][36]  = llr_new[4][7];
        llr_in_tmp[4][37]  = llr_new[4][8];
        llr_in_tmp[4][38]  = llr_new[4][9];
        llr_in_tmp[4][39]  = llr_new[4][10];
        llr_in_tmp[4][40]  = llr_new[4][11];
        llr_in_tmp[4][41]  = llr_new[4][12];
    end
 
    1:begin 
        llr_in_tmp[4][0]  = llr_new[4][27];
        llr_in_tmp[4][1]  = llr_new[4][28];
        llr_in_tmp[4][2]  = llr_new[4][29];
        llr_in_tmp[4][3]  = llr_new[4][30];
        llr_in_tmp[4][4]  = llr_new[4][31];
        llr_in_tmp[4][5]  = llr_new[4][32];
        llr_in_tmp[4][6]  = llr_new[4][33];
        llr_in_tmp[4][7]  = llr_new[4][34];
        llr_in_tmp[4][8]  = llr_new[4][35];
        llr_in_tmp[4][9]  = llr_new[4][36];
        llr_in_tmp[4][10]  = llr_new[4][37];
        llr_in_tmp[4][11]  = llr_new[4][38];
        llr_in_tmp[4][12]  = llr_new[4][39];
        llr_in_tmp[4][13]  = llr_new[4][40];
        llr_in_tmp[4][14]  = llr_new[4][41];
        llr_in_tmp[4][15]  = llr_new[4][0];
        llr_in_tmp[4][16]  = llr_new[4][1];
        llr_in_tmp[4][17]  = llr_new[4][2];
        llr_in_tmp[4][18]  = llr_new[4][3];
        llr_in_tmp[4][19]  = llr_new[4][4];
        llr_in_tmp[4][20]  = llr_new[4][5];
        llr_in_tmp[4][21]  = llr_new[4][6];
        llr_in_tmp[4][22]  = llr_new[4][7];
        llr_in_tmp[4][23]  = llr_new[4][8];
        llr_in_tmp[4][24]  = llr_new[4][9];
        llr_in_tmp[4][25]  = llr_new[4][10];
        llr_in_tmp[4][26]  = llr_new[4][11];
        llr_in_tmp[4][27]  = llr_new[4][12];
        llr_in_tmp[4][28]  = llr_new[4][13];
        llr_in_tmp[4][29]  = llr_new[4][14];
        llr_in_tmp[4][30]  = llr_new[4][15];
        llr_in_tmp[4][31]  = llr_new[4][16];
        llr_in_tmp[4][32]  = llr_new[4][17];
        llr_in_tmp[4][33]  = llr_new[4][18];
        llr_in_tmp[4][34]  = llr_new[4][19];
        llr_in_tmp[4][35]  = llr_new[4][20];
        llr_in_tmp[4][36]  = llr_new[4][21];
        llr_in_tmp[4][37]  = llr_new[4][22];
        llr_in_tmp[4][38]  = llr_new[4][23];
        llr_in_tmp[4][39]  = llr_new[4][24];
        llr_in_tmp[4][40]  = llr_new[4][25];
        llr_in_tmp[4][41]  = llr_new[4][26];
    end
 
    2:begin 
        llr_in_tmp[4][0]  = llr_new[4][0];
        llr_in_tmp[4][1]  = llr_new[4][1];
        llr_in_tmp[4][2]  = llr_new[4][2];
        llr_in_tmp[4][3]  = llr_new[4][3];
        llr_in_tmp[4][4]  = llr_new[4][4];
        llr_in_tmp[4][5]  = llr_new[4][5];
        llr_in_tmp[4][6]  = llr_new[4][6];
        llr_in_tmp[4][7]  = llr_new[4][7];
        llr_in_tmp[4][8]  = llr_new[4][8];
        llr_in_tmp[4][9]  = llr_new[4][9];
        llr_in_tmp[4][10]  = llr_new[4][10];
        llr_in_tmp[4][11]  = llr_new[4][11];
        llr_in_tmp[4][12]  = llr_new[4][12];
        llr_in_tmp[4][13]  = llr_new[4][13];
        llr_in_tmp[4][14]  = llr_new[4][14];
        llr_in_tmp[4][15]  = llr_new[4][15];
        llr_in_tmp[4][16]  = llr_new[4][16];
        llr_in_tmp[4][17]  = llr_new[4][17];
        llr_in_tmp[4][18]  = llr_new[4][18];
        llr_in_tmp[4][19]  = llr_new[4][19];
        llr_in_tmp[4][20]  = llr_new[4][20];
        llr_in_tmp[4][21]  = llr_new[4][21];
        llr_in_tmp[4][22]  = llr_new[4][22];
        llr_in_tmp[4][23]  = llr_new[4][23];
        llr_in_tmp[4][24]  = llr_new[4][24];
        llr_in_tmp[4][25]  = llr_new[4][25];
        llr_in_tmp[4][26]  = llr_new[4][26];
        llr_in_tmp[4][27]  = llr_new[4][27];
        llr_in_tmp[4][28]  = llr_new[4][28];
        llr_in_tmp[4][29]  = llr_new[4][29];
        llr_in_tmp[4][30]  = llr_new[4][30];
        llr_in_tmp[4][31]  = llr_new[4][31];
        llr_in_tmp[4][32]  = llr_new[4][32];
        llr_in_tmp[4][33]  = llr_new[4][33];
        llr_in_tmp[4][34]  = llr_new[4][34];
        llr_in_tmp[4][35]  = llr_new[4][35];
        llr_in_tmp[4][36]  = llr_new[4][36];
        llr_in_tmp[4][37]  = llr_new[4][37];
        llr_in_tmp[4][38]  = llr_new[4][38];
        llr_in_tmp[4][39]  = llr_new[4][39];
        llr_in_tmp[4][40]  = llr_new[4][40];
        llr_in_tmp[4][41]  = llr_new[4][41];
    end
 
    3:begin 
        llr_in_tmp[4][0]  = llr_new[4][0];
        llr_in_tmp[4][1]  = llr_new[4][1];
        llr_in_tmp[4][2]  = llr_new[4][2];
        llr_in_tmp[4][3]  = llr_new[4][3];
        llr_in_tmp[4][4]  = llr_new[4][4];
        llr_in_tmp[4][5]  = llr_new[4][5];
        llr_in_tmp[4][6]  = llr_new[4][6];
        llr_in_tmp[4][7]  = llr_new[4][7];
        llr_in_tmp[4][8]  = llr_new[4][8];
        llr_in_tmp[4][9]  = llr_new[4][9];
        llr_in_tmp[4][10]  = llr_new[4][10];
        llr_in_tmp[4][11]  = llr_new[4][11];
        llr_in_tmp[4][12]  = llr_new[4][12];
        llr_in_tmp[4][13]  = llr_new[4][13];
        llr_in_tmp[4][14]  = llr_new[4][14];
        llr_in_tmp[4][15]  = llr_new[4][15];
        llr_in_tmp[4][16]  = llr_new[4][16];
        llr_in_tmp[4][17]  = llr_new[4][17];
        llr_in_tmp[4][18]  = llr_new[4][18];
        llr_in_tmp[4][19]  = llr_new[4][19];
        llr_in_tmp[4][20]  = llr_new[4][20];
        llr_in_tmp[4][21]  = llr_new[4][21];
        llr_in_tmp[4][22]  = llr_new[4][22];
        llr_in_tmp[4][23]  = llr_new[4][23];
        llr_in_tmp[4][24]  = llr_new[4][24];
        llr_in_tmp[4][25]  = llr_new[4][25];
        llr_in_tmp[4][26]  = llr_new[4][26];
        llr_in_tmp[4][27]  = llr_new[4][27];
        llr_in_tmp[4][28]  = llr_new[4][28];
        llr_in_tmp[4][29]  = llr_new[4][29];
        llr_in_tmp[4][30]  = llr_new[4][30];
        llr_in_tmp[4][31]  = llr_new[4][31];
        llr_in_tmp[4][32]  = llr_new[4][32];
        llr_in_tmp[4][33]  = llr_new[4][33];
        llr_in_tmp[4][34]  = llr_new[4][34];
        llr_in_tmp[4][35]  = llr_new[4][35];
        llr_in_tmp[4][36]  = llr_new[4][36];
        llr_in_tmp[4][37]  = llr_new[4][37];
        llr_in_tmp[4][38]  = llr_new[4][38];
        llr_in_tmp[4][39]  = llr_new[4][39];
        llr_in_tmp[4][40]  = llr_new[4][40];
        llr_in_tmp[4][41]  = llr_new[4][41];
    end
 
    4:begin 
        llr_in_tmp[4][0]  = llr_new[4][40];
        llr_in_tmp[4][1]  = llr_new[4][41];
        llr_in_tmp[4][2]  = llr_new[4][0];
        llr_in_tmp[4][3]  = llr_new[4][1];
        llr_in_tmp[4][4]  = llr_new[4][2];
        llr_in_tmp[4][5]  = llr_new[4][3];
        llr_in_tmp[4][6]  = llr_new[4][4];
        llr_in_tmp[4][7]  = llr_new[4][5];
        llr_in_tmp[4][8]  = llr_new[4][6];
        llr_in_tmp[4][9]  = llr_new[4][7];
        llr_in_tmp[4][10]  = llr_new[4][8];
        llr_in_tmp[4][11]  = llr_new[4][9];
        llr_in_tmp[4][12]  = llr_new[4][10];
        llr_in_tmp[4][13]  = llr_new[4][11];
        llr_in_tmp[4][14]  = llr_new[4][12];
        llr_in_tmp[4][15]  = llr_new[4][13];
        llr_in_tmp[4][16]  = llr_new[4][14];
        llr_in_tmp[4][17]  = llr_new[4][15];
        llr_in_tmp[4][18]  = llr_new[4][16];
        llr_in_tmp[4][19]  = llr_new[4][17];
        llr_in_tmp[4][20]  = llr_new[4][18];
        llr_in_tmp[4][21]  = llr_new[4][19];
        llr_in_tmp[4][22]  = llr_new[4][20];
        llr_in_tmp[4][23]  = llr_new[4][21];
        llr_in_tmp[4][24]  = llr_new[4][22];
        llr_in_tmp[4][25]  = llr_new[4][23];
        llr_in_tmp[4][26]  = llr_new[4][24];
        llr_in_tmp[4][27]  = llr_new[4][25];
        llr_in_tmp[4][28]  = llr_new[4][26];
        llr_in_tmp[4][29]  = llr_new[4][27];
        llr_in_tmp[4][30]  = llr_new[4][28];
        llr_in_tmp[4][31]  = llr_new[4][29];
        llr_in_tmp[4][32]  = llr_new[4][30];
        llr_in_tmp[4][33]  = llr_new[4][31];
        llr_in_tmp[4][34]  = llr_new[4][32];
        llr_in_tmp[4][35]  = llr_new[4][33];
        llr_in_tmp[4][36]  = llr_new[4][34];
        llr_in_tmp[4][37]  = llr_new[4][35];
        llr_in_tmp[4][38]  = llr_new[4][36];
        llr_in_tmp[4][39]  = llr_new[4][37];
        llr_in_tmp[4][40]  = llr_new[4][38];
        llr_in_tmp[4][41]  = llr_new[4][39];
    end
 
    5:begin 
        llr_in_tmp[4][0]  = llr_new[4][0];
        llr_in_tmp[4][1]  = llr_new[4][1];
        llr_in_tmp[4][2]  = llr_new[4][2];
        llr_in_tmp[4][3]  = llr_new[4][3];
        llr_in_tmp[4][4]  = llr_new[4][4];
        llr_in_tmp[4][5]  = llr_new[4][5];
        llr_in_tmp[4][6]  = llr_new[4][6];
        llr_in_tmp[4][7]  = llr_new[4][7];
        llr_in_tmp[4][8]  = llr_new[4][8];
        llr_in_tmp[4][9]  = llr_new[4][9];
        llr_in_tmp[4][10]  = llr_new[4][10];
        llr_in_tmp[4][11]  = llr_new[4][11];
        llr_in_tmp[4][12]  = llr_new[4][12];
        llr_in_tmp[4][13]  = llr_new[4][13];
        llr_in_tmp[4][14]  = llr_new[4][14];
        llr_in_tmp[4][15]  = llr_new[4][15];
        llr_in_tmp[4][16]  = llr_new[4][16];
        llr_in_tmp[4][17]  = llr_new[4][17];
        llr_in_tmp[4][18]  = llr_new[4][18];
        llr_in_tmp[4][19]  = llr_new[4][19];
        llr_in_tmp[4][20]  = llr_new[4][20];
        llr_in_tmp[4][21]  = llr_new[4][21];
        llr_in_tmp[4][22]  = llr_new[4][22];
        llr_in_tmp[4][23]  = llr_new[4][23];
        llr_in_tmp[4][24]  = llr_new[4][24];
        llr_in_tmp[4][25]  = llr_new[4][25];
        llr_in_tmp[4][26]  = llr_new[4][26];
        llr_in_tmp[4][27]  = llr_new[4][27];
        llr_in_tmp[4][28]  = llr_new[4][28];
        llr_in_tmp[4][29]  = llr_new[4][29];
        llr_in_tmp[4][30]  = llr_new[4][30];
        llr_in_tmp[4][31]  = llr_new[4][31];
        llr_in_tmp[4][32]  = llr_new[4][32];
        llr_in_tmp[4][33]  = llr_new[4][33];
        llr_in_tmp[4][34]  = llr_new[4][34];
        llr_in_tmp[4][35]  = llr_new[4][35];
        llr_in_tmp[4][36]  = llr_new[4][36];
        llr_in_tmp[4][37]  = llr_new[4][37];
        llr_in_tmp[4][38]  = llr_new[4][38];
        llr_in_tmp[4][39]  = llr_new[4][39];
        llr_in_tmp[4][40]  = llr_new[4][40];
        llr_in_tmp[4][41]  = llr_new[4][41];
    end
 
    6:begin 
        llr_in_tmp[4][0]  = llr_new[4][0];
        llr_in_tmp[4][1]  = llr_new[4][1];
        llr_in_tmp[4][2]  = llr_new[4][2];
        llr_in_tmp[4][3]  = llr_new[4][3];
        llr_in_tmp[4][4]  = llr_new[4][4];
        llr_in_tmp[4][5]  = llr_new[4][5];
        llr_in_tmp[4][6]  = llr_new[4][6];
        llr_in_tmp[4][7]  = llr_new[4][7];
        llr_in_tmp[4][8]  = llr_new[4][8];
        llr_in_tmp[4][9]  = llr_new[4][9];
        llr_in_tmp[4][10]  = llr_new[4][10];
        llr_in_tmp[4][11]  = llr_new[4][11];
        llr_in_tmp[4][12]  = llr_new[4][12];
        llr_in_tmp[4][13]  = llr_new[4][13];
        llr_in_tmp[4][14]  = llr_new[4][14];
        llr_in_tmp[4][15]  = llr_new[4][15];
        llr_in_tmp[4][16]  = llr_new[4][16];
        llr_in_tmp[4][17]  = llr_new[4][17];
        llr_in_tmp[4][18]  = llr_new[4][18];
        llr_in_tmp[4][19]  = llr_new[4][19];
        llr_in_tmp[4][20]  = llr_new[4][20];
        llr_in_tmp[4][21]  = llr_new[4][21];
        llr_in_tmp[4][22]  = llr_new[4][22];
        llr_in_tmp[4][23]  = llr_new[4][23];
        llr_in_tmp[4][24]  = llr_new[4][24];
        llr_in_tmp[4][25]  = llr_new[4][25];
        llr_in_tmp[4][26]  = llr_new[4][26];
        llr_in_tmp[4][27]  = llr_new[4][27];
        llr_in_tmp[4][28]  = llr_new[4][28];
        llr_in_tmp[4][29]  = llr_new[4][29];
        llr_in_tmp[4][30]  = llr_new[4][30];
        llr_in_tmp[4][31]  = llr_new[4][31];
        llr_in_tmp[4][32]  = llr_new[4][32];
        llr_in_tmp[4][33]  = llr_new[4][33];
        llr_in_tmp[4][34]  = llr_new[4][34];
        llr_in_tmp[4][35]  = llr_new[4][35];
        llr_in_tmp[4][36]  = llr_new[4][36];
        llr_in_tmp[4][37]  = llr_new[4][37];
        llr_in_tmp[4][38]  = llr_new[4][38];
        llr_in_tmp[4][39]  = llr_new[4][39];
        llr_in_tmp[4][40]  = llr_new[4][40];
        llr_in_tmp[4][41]  = llr_new[4][41];
    end
 
    7:begin 
        llr_in_tmp[4][0]  = llr_new[4][31];
        llr_in_tmp[4][1]  = llr_new[4][32];
        llr_in_tmp[4][2]  = llr_new[4][33];
        llr_in_tmp[4][3]  = llr_new[4][34];
        llr_in_tmp[4][4]  = llr_new[4][35];
        llr_in_tmp[4][5]  = llr_new[4][36];
        llr_in_tmp[4][6]  = llr_new[4][37];
        llr_in_tmp[4][7]  = llr_new[4][38];
        llr_in_tmp[4][8]  = llr_new[4][39];
        llr_in_tmp[4][9]  = llr_new[4][40];
        llr_in_tmp[4][10]  = llr_new[4][41];
        llr_in_tmp[4][11]  = llr_new[4][0];
        llr_in_tmp[4][12]  = llr_new[4][1];
        llr_in_tmp[4][13]  = llr_new[4][2];
        llr_in_tmp[4][14]  = llr_new[4][3];
        llr_in_tmp[4][15]  = llr_new[4][4];
        llr_in_tmp[4][16]  = llr_new[4][5];
        llr_in_tmp[4][17]  = llr_new[4][6];
        llr_in_tmp[4][18]  = llr_new[4][7];
        llr_in_tmp[4][19]  = llr_new[4][8];
        llr_in_tmp[4][20]  = llr_new[4][9];
        llr_in_tmp[4][21]  = llr_new[4][10];
        llr_in_tmp[4][22]  = llr_new[4][11];
        llr_in_tmp[4][23]  = llr_new[4][12];
        llr_in_tmp[4][24]  = llr_new[4][13];
        llr_in_tmp[4][25]  = llr_new[4][14];
        llr_in_tmp[4][26]  = llr_new[4][15];
        llr_in_tmp[4][27]  = llr_new[4][16];
        llr_in_tmp[4][28]  = llr_new[4][17];
        llr_in_tmp[4][29]  = llr_new[4][18];
        llr_in_tmp[4][30]  = llr_new[4][19];
        llr_in_tmp[4][31]  = llr_new[4][20];
        llr_in_tmp[4][32]  = llr_new[4][21];
        llr_in_tmp[4][33]  = llr_new[4][22];
        llr_in_tmp[4][34]  = llr_new[4][23];
        llr_in_tmp[4][35]  = llr_new[4][24];
        llr_in_tmp[4][36]  = llr_new[4][25];
        llr_in_tmp[4][37]  = llr_new[4][26];
        llr_in_tmp[4][38]  = llr_new[4][27];
        llr_in_tmp[4][39]  = llr_new[4][28];
        llr_in_tmp[4][40]  = llr_new[4][29];
        llr_in_tmp[4][41]  = llr_new[4][30];
    end
 
endcase
end

if (chk_n_input_valid) begin
case (curr_layer)
    0:begin 
        llr_in_tmp[5][0]  = llr_new[5][0];
        llr_in_tmp[5][1]  = llr_new[5][1];
        llr_in_tmp[5][2]  = llr_new[5][2];
        llr_in_tmp[5][3]  = llr_new[5][3];
        llr_in_tmp[5][4]  = llr_new[5][4];
        llr_in_tmp[5][5]  = llr_new[5][5];
        llr_in_tmp[5][6]  = llr_new[5][6];
        llr_in_tmp[5][7]  = llr_new[5][7];
        llr_in_tmp[5][8]  = llr_new[5][8];
        llr_in_tmp[5][9]  = llr_new[5][9];
        llr_in_tmp[5][10]  = llr_new[5][10];
        llr_in_tmp[5][11]  = llr_new[5][11];
        llr_in_tmp[5][12]  = llr_new[5][12];
        llr_in_tmp[5][13]  = llr_new[5][13];
        llr_in_tmp[5][14]  = llr_new[5][14];
        llr_in_tmp[5][15]  = llr_new[5][15];
        llr_in_tmp[5][16]  = llr_new[5][16];
        llr_in_tmp[5][17]  = llr_new[5][17];
        llr_in_tmp[5][18]  = llr_new[5][18];
        llr_in_tmp[5][19]  = llr_new[5][19];
        llr_in_tmp[5][20]  = llr_new[5][20];
        llr_in_tmp[5][21]  = llr_new[5][21];
        llr_in_tmp[5][22]  = llr_new[5][22];
        llr_in_tmp[5][23]  = llr_new[5][23];
        llr_in_tmp[5][24]  = llr_new[5][24];
        llr_in_tmp[5][25]  = llr_new[5][25];
        llr_in_tmp[5][26]  = llr_new[5][26];
        llr_in_tmp[5][27]  = llr_new[5][27];
        llr_in_tmp[5][28]  = llr_new[5][28];
        llr_in_tmp[5][29]  = llr_new[5][29];
        llr_in_tmp[5][30]  = llr_new[5][30];
        llr_in_tmp[5][31]  = llr_new[5][31];
        llr_in_tmp[5][32]  = llr_new[5][32];
        llr_in_tmp[5][33]  = llr_new[5][33];
        llr_in_tmp[5][34]  = llr_new[5][34];
        llr_in_tmp[5][35]  = llr_new[5][35];
        llr_in_tmp[5][36]  = llr_new[5][36];
        llr_in_tmp[5][37]  = llr_new[5][37];
        llr_in_tmp[5][38]  = llr_new[5][38];
        llr_in_tmp[5][39]  = llr_new[5][39];
        llr_in_tmp[5][40]  = llr_new[5][40];
        llr_in_tmp[5][41]  = llr_new[5][41];
    end
 
    1:begin 
        llr_in_tmp[5][0]  = llr_new[5][0];
        llr_in_tmp[5][1]  = llr_new[5][1];
        llr_in_tmp[5][2]  = llr_new[5][2];
        llr_in_tmp[5][3]  = llr_new[5][3];
        llr_in_tmp[5][4]  = llr_new[5][4];
        llr_in_tmp[5][5]  = llr_new[5][5];
        llr_in_tmp[5][6]  = llr_new[5][6];
        llr_in_tmp[5][7]  = llr_new[5][7];
        llr_in_tmp[5][8]  = llr_new[5][8];
        llr_in_tmp[5][9]  = llr_new[5][9];
        llr_in_tmp[5][10]  = llr_new[5][10];
        llr_in_tmp[5][11]  = llr_new[5][11];
        llr_in_tmp[5][12]  = llr_new[5][12];
        llr_in_tmp[5][13]  = llr_new[5][13];
        llr_in_tmp[5][14]  = llr_new[5][14];
        llr_in_tmp[5][15]  = llr_new[5][15];
        llr_in_tmp[5][16]  = llr_new[5][16];
        llr_in_tmp[5][17]  = llr_new[5][17];
        llr_in_tmp[5][18]  = llr_new[5][18];
        llr_in_tmp[5][19]  = llr_new[5][19];
        llr_in_tmp[5][20]  = llr_new[5][20];
        llr_in_tmp[5][21]  = llr_new[5][21];
        llr_in_tmp[5][22]  = llr_new[5][22];
        llr_in_tmp[5][23]  = llr_new[5][23];
        llr_in_tmp[5][24]  = llr_new[5][24];
        llr_in_tmp[5][25]  = llr_new[5][25];
        llr_in_tmp[5][26]  = llr_new[5][26];
        llr_in_tmp[5][27]  = llr_new[5][27];
        llr_in_tmp[5][28]  = llr_new[5][28];
        llr_in_tmp[5][29]  = llr_new[5][29];
        llr_in_tmp[5][30]  = llr_new[5][30];
        llr_in_tmp[5][31]  = llr_new[5][31];
        llr_in_tmp[5][32]  = llr_new[5][32];
        llr_in_tmp[5][33]  = llr_new[5][33];
        llr_in_tmp[5][34]  = llr_new[5][34];
        llr_in_tmp[5][35]  = llr_new[5][35];
        llr_in_tmp[5][36]  = llr_new[5][36];
        llr_in_tmp[5][37]  = llr_new[5][37];
        llr_in_tmp[5][38]  = llr_new[5][38];
        llr_in_tmp[5][39]  = llr_new[5][39];
        llr_in_tmp[5][40]  = llr_new[5][40];
        llr_in_tmp[5][41]  = llr_new[5][41];
    end
 
    2:begin 
        llr_in_tmp[5][0]  = llr_new[5][7];
        llr_in_tmp[5][1]  = llr_new[5][8];
        llr_in_tmp[5][2]  = llr_new[5][9];
        llr_in_tmp[5][3]  = llr_new[5][10];
        llr_in_tmp[5][4]  = llr_new[5][11];
        llr_in_tmp[5][5]  = llr_new[5][12];
        llr_in_tmp[5][6]  = llr_new[5][13];
        llr_in_tmp[5][7]  = llr_new[5][14];
        llr_in_tmp[5][8]  = llr_new[5][15];
        llr_in_tmp[5][9]  = llr_new[5][16];
        llr_in_tmp[5][10]  = llr_new[5][17];
        llr_in_tmp[5][11]  = llr_new[5][18];
        llr_in_tmp[5][12]  = llr_new[5][19];
        llr_in_tmp[5][13]  = llr_new[5][20];
        llr_in_tmp[5][14]  = llr_new[5][21];
        llr_in_tmp[5][15]  = llr_new[5][22];
        llr_in_tmp[5][16]  = llr_new[5][23];
        llr_in_tmp[5][17]  = llr_new[5][24];
        llr_in_tmp[5][18]  = llr_new[5][25];
        llr_in_tmp[5][19]  = llr_new[5][26];
        llr_in_tmp[5][20]  = llr_new[5][27];
        llr_in_tmp[5][21]  = llr_new[5][28];
        llr_in_tmp[5][22]  = llr_new[5][29];
        llr_in_tmp[5][23]  = llr_new[5][30];
        llr_in_tmp[5][24]  = llr_new[5][31];
        llr_in_tmp[5][25]  = llr_new[5][32];
        llr_in_tmp[5][26]  = llr_new[5][33];
        llr_in_tmp[5][27]  = llr_new[5][34];
        llr_in_tmp[5][28]  = llr_new[5][35];
        llr_in_tmp[5][29]  = llr_new[5][36];
        llr_in_tmp[5][30]  = llr_new[5][37];
        llr_in_tmp[5][31]  = llr_new[5][38];
        llr_in_tmp[5][32]  = llr_new[5][39];
        llr_in_tmp[5][33]  = llr_new[5][40];
        llr_in_tmp[5][34]  = llr_new[5][41];
        llr_in_tmp[5][35]  = llr_new[5][0];
        llr_in_tmp[5][36]  = llr_new[5][1];
        llr_in_tmp[5][37]  = llr_new[5][2];
        llr_in_tmp[5][38]  = llr_new[5][3];
        llr_in_tmp[5][39]  = llr_new[5][4];
        llr_in_tmp[5][40]  = llr_new[5][5];
        llr_in_tmp[5][41]  = llr_new[5][6];
    end
 
    3:begin 
        llr_in_tmp[5][0]  = llr_new[5][12];
        llr_in_tmp[5][1]  = llr_new[5][13];
        llr_in_tmp[5][2]  = llr_new[5][14];
        llr_in_tmp[5][3]  = llr_new[5][15];
        llr_in_tmp[5][4]  = llr_new[5][16];
        llr_in_tmp[5][5]  = llr_new[5][17];
        llr_in_tmp[5][6]  = llr_new[5][18];
        llr_in_tmp[5][7]  = llr_new[5][19];
        llr_in_tmp[5][8]  = llr_new[5][20];
        llr_in_tmp[5][9]  = llr_new[5][21];
        llr_in_tmp[5][10]  = llr_new[5][22];
        llr_in_tmp[5][11]  = llr_new[5][23];
        llr_in_tmp[5][12]  = llr_new[5][24];
        llr_in_tmp[5][13]  = llr_new[5][25];
        llr_in_tmp[5][14]  = llr_new[5][26];
        llr_in_tmp[5][15]  = llr_new[5][27];
        llr_in_tmp[5][16]  = llr_new[5][28];
        llr_in_tmp[5][17]  = llr_new[5][29];
        llr_in_tmp[5][18]  = llr_new[5][30];
        llr_in_tmp[5][19]  = llr_new[5][31];
        llr_in_tmp[5][20]  = llr_new[5][32];
        llr_in_tmp[5][21]  = llr_new[5][33];
        llr_in_tmp[5][22]  = llr_new[5][34];
        llr_in_tmp[5][23]  = llr_new[5][35];
        llr_in_tmp[5][24]  = llr_new[5][36];
        llr_in_tmp[5][25]  = llr_new[5][37];
        llr_in_tmp[5][26]  = llr_new[5][38];
        llr_in_tmp[5][27]  = llr_new[5][39];
        llr_in_tmp[5][28]  = llr_new[5][40];
        llr_in_tmp[5][29]  = llr_new[5][41];
        llr_in_tmp[5][30]  = llr_new[5][0];
        llr_in_tmp[5][31]  = llr_new[5][1];
        llr_in_tmp[5][32]  = llr_new[5][2];
        llr_in_tmp[5][33]  = llr_new[5][3];
        llr_in_tmp[5][34]  = llr_new[5][4];
        llr_in_tmp[5][35]  = llr_new[5][5];
        llr_in_tmp[5][36]  = llr_new[5][6];
        llr_in_tmp[5][37]  = llr_new[5][7];
        llr_in_tmp[5][38]  = llr_new[5][8];
        llr_in_tmp[5][39]  = llr_new[5][9];
        llr_in_tmp[5][40]  = llr_new[5][10];
        llr_in_tmp[5][41]  = llr_new[5][11];
    end
 
    4:begin 
        llr_in_tmp[5][0]  = llr_new[5][0];
        llr_in_tmp[5][1]  = llr_new[5][1];
        llr_in_tmp[5][2]  = llr_new[5][2];
        llr_in_tmp[5][3]  = llr_new[5][3];
        llr_in_tmp[5][4]  = llr_new[5][4];
        llr_in_tmp[5][5]  = llr_new[5][5];
        llr_in_tmp[5][6]  = llr_new[5][6];
        llr_in_tmp[5][7]  = llr_new[5][7];
        llr_in_tmp[5][8]  = llr_new[5][8];
        llr_in_tmp[5][9]  = llr_new[5][9];
        llr_in_tmp[5][10]  = llr_new[5][10];
        llr_in_tmp[5][11]  = llr_new[5][11];
        llr_in_tmp[5][12]  = llr_new[5][12];
        llr_in_tmp[5][13]  = llr_new[5][13];
        llr_in_tmp[5][14]  = llr_new[5][14];
        llr_in_tmp[5][15]  = llr_new[5][15];
        llr_in_tmp[5][16]  = llr_new[5][16];
        llr_in_tmp[5][17]  = llr_new[5][17];
        llr_in_tmp[5][18]  = llr_new[5][18];
        llr_in_tmp[5][19]  = llr_new[5][19];
        llr_in_tmp[5][20]  = llr_new[5][20];
        llr_in_tmp[5][21]  = llr_new[5][21];
        llr_in_tmp[5][22]  = llr_new[5][22];
        llr_in_tmp[5][23]  = llr_new[5][23];
        llr_in_tmp[5][24]  = llr_new[5][24];
        llr_in_tmp[5][25]  = llr_new[5][25];
        llr_in_tmp[5][26]  = llr_new[5][26];
        llr_in_tmp[5][27]  = llr_new[5][27];
        llr_in_tmp[5][28]  = llr_new[5][28];
        llr_in_tmp[5][29]  = llr_new[5][29];
        llr_in_tmp[5][30]  = llr_new[5][30];
        llr_in_tmp[5][31]  = llr_new[5][31];
        llr_in_tmp[5][32]  = llr_new[5][32];
        llr_in_tmp[5][33]  = llr_new[5][33];
        llr_in_tmp[5][34]  = llr_new[5][34];
        llr_in_tmp[5][35]  = llr_new[5][35];
        llr_in_tmp[5][36]  = llr_new[5][36];
        llr_in_tmp[5][37]  = llr_new[5][37];
        llr_in_tmp[5][38]  = llr_new[5][38];
        llr_in_tmp[5][39]  = llr_new[5][39];
        llr_in_tmp[5][40]  = llr_new[5][40];
        llr_in_tmp[5][41]  = llr_new[5][41];
    end
 
    5:begin 
        llr_in_tmp[5][0]  = llr_new[5][22];
        llr_in_tmp[5][1]  = llr_new[5][23];
        llr_in_tmp[5][2]  = llr_new[5][24];
        llr_in_tmp[5][3]  = llr_new[5][25];
        llr_in_tmp[5][4]  = llr_new[5][26];
        llr_in_tmp[5][5]  = llr_new[5][27];
        llr_in_tmp[5][6]  = llr_new[5][28];
        llr_in_tmp[5][7]  = llr_new[5][29];
        llr_in_tmp[5][8]  = llr_new[5][30];
        llr_in_tmp[5][9]  = llr_new[5][31];
        llr_in_tmp[5][10]  = llr_new[5][32];
        llr_in_tmp[5][11]  = llr_new[5][33];
        llr_in_tmp[5][12]  = llr_new[5][34];
        llr_in_tmp[5][13]  = llr_new[5][35];
        llr_in_tmp[5][14]  = llr_new[5][36];
        llr_in_tmp[5][15]  = llr_new[5][37];
        llr_in_tmp[5][16]  = llr_new[5][38];
        llr_in_tmp[5][17]  = llr_new[5][39];
        llr_in_tmp[5][18]  = llr_new[5][40];
        llr_in_tmp[5][19]  = llr_new[5][41];
        llr_in_tmp[5][20]  = llr_new[5][0];
        llr_in_tmp[5][21]  = llr_new[5][1];
        llr_in_tmp[5][22]  = llr_new[5][2];
        llr_in_tmp[5][23]  = llr_new[5][3];
        llr_in_tmp[5][24]  = llr_new[5][4];
        llr_in_tmp[5][25]  = llr_new[5][5];
        llr_in_tmp[5][26]  = llr_new[5][6];
        llr_in_tmp[5][27]  = llr_new[5][7];
        llr_in_tmp[5][28]  = llr_new[5][8];
        llr_in_tmp[5][29]  = llr_new[5][9];
        llr_in_tmp[5][30]  = llr_new[5][10];
        llr_in_tmp[5][31]  = llr_new[5][11];
        llr_in_tmp[5][32]  = llr_new[5][12];
        llr_in_tmp[5][33]  = llr_new[5][13];
        llr_in_tmp[5][34]  = llr_new[5][14];
        llr_in_tmp[5][35]  = llr_new[5][15];
        llr_in_tmp[5][36]  = llr_new[5][16];
        llr_in_tmp[5][37]  = llr_new[5][17];
        llr_in_tmp[5][38]  = llr_new[5][18];
        llr_in_tmp[5][39]  = llr_new[5][19];
        llr_in_tmp[5][40]  = llr_new[5][20];
        llr_in_tmp[5][41]  = llr_new[5][21];
    end
 
    6:begin 
        llr_in_tmp[5][0]  = llr_new[5][21];
        llr_in_tmp[5][1]  = llr_new[5][22];
        llr_in_tmp[5][2]  = llr_new[5][23];
        llr_in_tmp[5][3]  = llr_new[5][24];
        llr_in_tmp[5][4]  = llr_new[5][25];
        llr_in_tmp[5][5]  = llr_new[5][26];
        llr_in_tmp[5][6]  = llr_new[5][27];
        llr_in_tmp[5][7]  = llr_new[5][28];
        llr_in_tmp[5][8]  = llr_new[5][29];
        llr_in_tmp[5][9]  = llr_new[5][30];
        llr_in_tmp[5][10]  = llr_new[5][31];
        llr_in_tmp[5][11]  = llr_new[5][32];
        llr_in_tmp[5][12]  = llr_new[5][33];
        llr_in_tmp[5][13]  = llr_new[5][34];
        llr_in_tmp[5][14]  = llr_new[5][35];
        llr_in_tmp[5][15]  = llr_new[5][36];
        llr_in_tmp[5][16]  = llr_new[5][37];
        llr_in_tmp[5][17]  = llr_new[5][38];
        llr_in_tmp[5][18]  = llr_new[5][39];
        llr_in_tmp[5][19]  = llr_new[5][40];
        llr_in_tmp[5][20]  = llr_new[5][41];
        llr_in_tmp[5][21]  = llr_new[5][0];
        llr_in_tmp[5][22]  = llr_new[5][1];
        llr_in_tmp[5][23]  = llr_new[5][2];
        llr_in_tmp[5][24]  = llr_new[5][3];
        llr_in_tmp[5][25]  = llr_new[5][4];
        llr_in_tmp[5][26]  = llr_new[5][5];
        llr_in_tmp[5][27]  = llr_new[5][6];
        llr_in_tmp[5][28]  = llr_new[5][7];
        llr_in_tmp[5][29]  = llr_new[5][8];
        llr_in_tmp[5][30]  = llr_new[5][9];
        llr_in_tmp[5][31]  = llr_new[5][10];
        llr_in_tmp[5][32]  = llr_new[5][11];
        llr_in_tmp[5][33]  = llr_new[5][12];
        llr_in_tmp[5][34]  = llr_new[5][13];
        llr_in_tmp[5][35]  = llr_new[5][14];
        llr_in_tmp[5][36]  = llr_new[5][15];
        llr_in_tmp[5][37]  = llr_new[5][16];
        llr_in_tmp[5][38]  = llr_new[5][17];
        llr_in_tmp[5][39]  = llr_new[5][18];
        llr_in_tmp[5][40]  = llr_new[5][19];
        llr_in_tmp[5][41]  = llr_new[5][20];
    end
 
    7:begin 
        llr_in_tmp[5][0]  = llr_new[5][0];
        llr_in_tmp[5][1]  = llr_new[5][1];
        llr_in_tmp[5][2]  = llr_new[5][2];
        llr_in_tmp[5][3]  = llr_new[5][3];
        llr_in_tmp[5][4]  = llr_new[5][4];
        llr_in_tmp[5][5]  = llr_new[5][5];
        llr_in_tmp[5][6]  = llr_new[5][6];
        llr_in_tmp[5][7]  = llr_new[5][7];
        llr_in_tmp[5][8]  = llr_new[5][8];
        llr_in_tmp[5][9]  = llr_new[5][9];
        llr_in_tmp[5][10]  = llr_new[5][10];
        llr_in_tmp[5][11]  = llr_new[5][11];
        llr_in_tmp[5][12]  = llr_new[5][12];
        llr_in_tmp[5][13]  = llr_new[5][13];
        llr_in_tmp[5][14]  = llr_new[5][14];
        llr_in_tmp[5][15]  = llr_new[5][15];
        llr_in_tmp[5][16]  = llr_new[5][16];
        llr_in_tmp[5][17]  = llr_new[5][17];
        llr_in_tmp[5][18]  = llr_new[5][18];
        llr_in_tmp[5][19]  = llr_new[5][19];
        llr_in_tmp[5][20]  = llr_new[5][20];
        llr_in_tmp[5][21]  = llr_new[5][21];
        llr_in_tmp[5][22]  = llr_new[5][22];
        llr_in_tmp[5][23]  = llr_new[5][23];
        llr_in_tmp[5][24]  = llr_new[5][24];
        llr_in_tmp[5][25]  = llr_new[5][25];
        llr_in_tmp[5][26]  = llr_new[5][26];
        llr_in_tmp[5][27]  = llr_new[5][27];
        llr_in_tmp[5][28]  = llr_new[5][28];
        llr_in_tmp[5][29]  = llr_new[5][29];
        llr_in_tmp[5][30]  = llr_new[5][30];
        llr_in_tmp[5][31]  = llr_new[5][31];
        llr_in_tmp[5][32]  = llr_new[5][32];
        llr_in_tmp[5][33]  = llr_new[5][33];
        llr_in_tmp[5][34]  = llr_new[5][34];
        llr_in_tmp[5][35]  = llr_new[5][35];
        llr_in_tmp[5][36]  = llr_new[5][36];
        llr_in_tmp[5][37]  = llr_new[5][37];
        llr_in_tmp[5][38]  = llr_new[5][38];
        llr_in_tmp[5][39]  = llr_new[5][39];
        llr_in_tmp[5][40]  = llr_new[5][40];
        llr_in_tmp[5][41]  = llr_new[5][41];
    end
 
endcase
end

if (chk_n_input_valid) begin
case (curr_layer)
    0:begin 
        llr_in_tmp[6][0]  = llr_new[6][5];
        llr_in_tmp[6][1]  = llr_new[6][6];
        llr_in_tmp[6][2]  = llr_new[6][7];
        llr_in_tmp[6][3]  = llr_new[6][8];
        llr_in_tmp[6][4]  = llr_new[6][9];
        llr_in_tmp[6][5]  = llr_new[6][10];
        llr_in_tmp[6][6]  = llr_new[6][11];
        llr_in_tmp[6][7]  = llr_new[6][12];
        llr_in_tmp[6][8]  = llr_new[6][13];
        llr_in_tmp[6][9]  = llr_new[6][14];
        llr_in_tmp[6][10]  = llr_new[6][15];
        llr_in_tmp[6][11]  = llr_new[6][16];
        llr_in_tmp[6][12]  = llr_new[6][17];
        llr_in_tmp[6][13]  = llr_new[6][18];
        llr_in_tmp[6][14]  = llr_new[6][19];
        llr_in_tmp[6][15]  = llr_new[6][20];
        llr_in_tmp[6][16]  = llr_new[6][21];
        llr_in_tmp[6][17]  = llr_new[6][22];
        llr_in_tmp[6][18]  = llr_new[6][23];
        llr_in_tmp[6][19]  = llr_new[6][24];
        llr_in_tmp[6][20]  = llr_new[6][25];
        llr_in_tmp[6][21]  = llr_new[6][26];
        llr_in_tmp[6][22]  = llr_new[6][27];
        llr_in_tmp[6][23]  = llr_new[6][28];
        llr_in_tmp[6][24]  = llr_new[6][29];
        llr_in_tmp[6][25]  = llr_new[6][30];
        llr_in_tmp[6][26]  = llr_new[6][31];
        llr_in_tmp[6][27]  = llr_new[6][32];
        llr_in_tmp[6][28]  = llr_new[6][33];
        llr_in_tmp[6][29]  = llr_new[6][34];
        llr_in_tmp[6][30]  = llr_new[6][35];
        llr_in_tmp[6][31]  = llr_new[6][36];
        llr_in_tmp[6][32]  = llr_new[6][37];
        llr_in_tmp[6][33]  = llr_new[6][38];
        llr_in_tmp[6][34]  = llr_new[6][39];
        llr_in_tmp[6][35]  = llr_new[6][40];
        llr_in_tmp[6][36]  = llr_new[6][41];
        llr_in_tmp[6][37]  = llr_new[6][0];
        llr_in_tmp[6][38]  = llr_new[6][1];
        llr_in_tmp[6][39]  = llr_new[6][2];
        llr_in_tmp[6][40]  = llr_new[6][3];
        llr_in_tmp[6][41]  = llr_new[6][4];
    end
 
    1:begin 
        llr_in_tmp[6][0]  = llr_new[6][0];
        llr_in_tmp[6][1]  = llr_new[6][1];
        llr_in_tmp[6][2]  = llr_new[6][2];
        llr_in_tmp[6][3]  = llr_new[6][3];
        llr_in_tmp[6][4]  = llr_new[6][4];
        llr_in_tmp[6][5]  = llr_new[6][5];
        llr_in_tmp[6][6]  = llr_new[6][6];
        llr_in_tmp[6][7]  = llr_new[6][7];
        llr_in_tmp[6][8]  = llr_new[6][8];
        llr_in_tmp[6][9]  = llr_new[6][9];
        llr_in_tmp[6][10]  = llr_new[6][10];
        llr_in_tmp[6][11]  = llr_new[6][11];
        llr_in_tmp[6][12]  = llr_new[6][12];
        llr_in_tmp[6][13]  = llr_new[6][13];
        llr_in_tmp[6][14]  = llr_new[6][14];
        llr_in_tmp[6][15]  = llr_new[6][15];
        llr_in_tmp[6][16]  = llr_new[6][16];
        llr_in_tmp[6][17]  = llr_new[6][17];
        llr_in_tmp[6][18]  = llr_new[6][18];
        llr_in_tmp[6][19]  = llr_new[6][19];
        llr_in_tmp[6][20]  = llr_new[6][20];
        llr_in_tmp[6][21]  = llr_new[6][21];
        llr_in_tmp[6][22]  = llr_new[6][22];
        llr_in_tmp[6][23]  = llr_new[6][23];
        llr_in_tmp[6][24]  = llr_new[6][24];
        llr_in_tmp[6][25]  = llr_new[6][25];
        llr_in_tmp[6][26]  = llr_new[6][26];
        llr_in_tmp[6][27]  = llr_new[6][27];
        llr_in_tmp[6][28]  = llr_new[6][28];
        llr_in_tmp[6][29]  = llr_new[6][29];
        llr_in_tmp[6][30]  = llr_new[6][30];
        llr_in_tmp[6][31]  = llr_new[6][31];
        llr_in_tmp[6][32]  = llr_new[6][32];
        llr_in_tmp[6][33]  = llr_new[6][33];
        llr_in_tmp[6][34]  = llr_new[6][34];
        llr_in_tmp[6][35]  = llr_new[6][35];
        llr_in_tmp[6][36]  = llr_new[6][36];
        llr_in_tmp[6][37]  = llr_new[6][37];
        llr_in_tmp[6][38]  = llr_new[6][38];
        llr_in_tmp[6][39]  = llr_new[6][39];
        llr_in_tmp[6][40]  = llr_new[6][40];
        llr_in_tmp[6][41]  = llr_new[6][41];
    end
 
    2:begin 
        llr_in_tmp[6][0]  = llr_new[6][0];
        llr_in_tmp[6][1]  = llr_new[6][1];
        llr_in_tmp[6][2]  = llr_new[6][2];
        llr_in_tmp[6][3]  = llr_new[6][3];
        llr_in_tmp[6][4]  = llr_new[6][4];
        llr_in_tmp[6][5]  = llr_new[6][5];
        llr_in_tmp[6][6]  = llr_new[6][6];
        llr_in_tmp[6][7]  = llr_new[6][7];
        llr_in_tmp[6][8]  = llr_new[6][8];
        llr_in_tmp[6][9]  = llr_new[6][9];
        llr_in_tmp[6][10]  = llr_new[6][10];
        llr_in_tmp[6][11]  = llr_new[6][11];
        llr_in_tmp[6][12]  = llr_new[6][12];
        llr_in_tmp[6][13]  = llr_new[6][13];
        llr_in_tmp[6][14]  = llr_new[6][14];
        llr_in_tmp[6][15]  = llr_new[6][15];
        llr_in_tmp[6][16]  = llr_new[6][16];
        llr_in_tmp[6][17]  = llr_new[6][17];
        llr_in_tmp[6][18]  = llr_new[6][18];
        llr_in_tmp[6][19]  = llr_new[6][19];
        llr_in_tmp[6][20]  = llr_new[6][20];
        llr_in_tmp[6][21]  = llr_new[6][21];
        llr_in_tmp[6][22]  = llr_new[6][22];
        llr_in_tmp[6][23]  = llr_new[6][23];
        llr_in_tmp[6][24]  = llr_new[6][24];
        llr_in_tmp[6][25]  = llr_new[6][25];
        llr_in_tmp[6][26]  = llr_new[6][26];
        llr_in_tmp[6][27]  = llr_new[6][27];
        llr_in_tmp[6][28]  = llr_new[6][28];
        llr_in_tmp[6][29]  = llr_new[6][29];
        llr_in_tmp[6][30]  = llr_new[6][30];
        llr_in_tmp[6][31]  = llr_new[6][31];
        llr_in_tmp[6][32]  = llr_new[6][32];
        llr_in_tmp[6][33]  = llr_new[6][33];
        llr_in_tmp[6][34]  = llr_new[6][34];
        llr_in_tmp[6][35]  = llr_new[6][35];
        llr_in_tmp[6][36]  = llr_new[6][36];
        llr_in_tmp[6][37]  = llr_new[6][37];
        llr_in_tmp[6][38]  = llr_new[6][38];
        llr_in_tmp[6][39]  = llr_new[6][39];
        llr_in_tmp[6][40]  = llr_new[6][40];
        llr_in_tmp[6][41]  = llr_new[6][41];
    end
 
    3:begin 
        llr_in_tmp[6][0]  = llr_new[6][20];
        llr_in_tmp[6][1]  = llr_new[6][21];
        llr_in_tmp[6][2]  = llr_new[6][22];
        llr_in_tmp[6][3]  = llr_new[6][23];
        llr_in_tmp[6][4]  = llr_new[6][24];
        llr_in_tmp[6][5]  = llr_new[6][25];
        llr_in_tmp[6][6]  = llr_new[6][26];
        llr_in_tmp[6][7]  = llr_new[6][27];
        llr_in_tmp[6][8]  = llr_new[6][28];
        llr_in_tmp[6][9]  = llr_new[6][29];
        llr_in_tmp[6][10]  = llr_new[6][30];
        llr_in_tmp[6][11]  = llr_new[6][31];
        llr_in_tmp[6][12]  = llr_new[6][32];
        llr_in_tmp[6][13]  = llr_new[6][33];
        llr_in_tmp[6][14]  = llr_new[6][34];
        llr_in_tmp[6][15]  = llr_new[6][35];
        llr_in_tmp[6][16]  = llr_new[6][36];
        llr_in_tmp[6][17]  = llr_new[6][37];
        llr_in_tmp[6][18]  = llr_new[6][38];
        llr_in_tmp[6][19]  = llr_new[6][39];
        llr_in_tmp[6][20]  = llr_new[6][40];
        llr_in_tmp[6][21]  = llr_new[6][41];
        llr_in_tmp[6][22]  = llr_new[6][0];
        llr_in_tmp[6][23]  = llr_new[6][1];
        llr_in_tmp[6][24]  = llr_new[6][2];
        llr_in_tmp[6][25]  = llr_new[6][3];
        llr_in_tmp[6][26]  = llr_new[6][4];
        llr_in_tmp[6][27]  = llr_new[6][5];
        llr_in_tmp[6][28]  = llr_new[6][6];
        llr_in_tmp[6][29]  = llr_new[6][7];
        llr_in_tmp[6][30]  = llr_new[6][8];
        llr_in_tmp[6][31]  = llr_new[6][9];
        llr_in_tmp[6][32]  = llr_new[6][10];
        llr_in_tmp[6][33]  = llr_new[6][11];
        llr_in_tmp[6][34]  = llr_new[6][12];
        llr_in_tmp[6][35]  = llr_new[6][13];
        llr_in_tmp[6][36]  = llr_new[6][14];
        llr_in_tmp[6][37]  = llr_new[6][15];
        llr_in_tmp[6][38]  = llr_new[6][16];
        llr_in_tmp[6][39]  = llr_new[6][17];
        llr_in_tmp[6][40]  = llr_new[6][18];
        llr_in_tmp[6][41]  = llr_new[6][19];
    end
 
    4:begin 
        llr_in_tmp[6][0]  = llr_new[6][39];
        llr_in_tmp[6][1]  = llr_new[6][40];
        llr_in_tmp[6][2]  = llr_new[6][41];
        llr_in_tmp[6][3]  = llr_new[6][0];
        llr_in_tmp[6][4]  = llr_new[6][1];
        llr_in_tmp[6][5]  = llr_new[6][2];
        llr_in_tmp[6][6]  = llr_new[6][3];
        llr_in_tmp[6][7]  = llr_new[6][4];
        llr_in_tmp[6][8]  = llr_new[6][5];
        llr_in_tmp[6][9]  = llr_new[6][6];
        llr_in_tmp[6][10]  = llr_new[6][7];
        llr_in_tmp[6][11]  = llr_new[6][8];
        llr_in_tmp[6][12]  = llr_new[6][9];
        llr_in_tmp[6][13]  = llr_new[6][10];
        llr_in_tmp[6][14]  = llr_new[6][11];
        llr_in_tmp[6][15]  = llr_new[6][12];
        llr_in_tmp[6][16]  = llr_new[6][13];
        llr_in_tmp[6][17]  = llr_new[6][14];
        llr_in_tmp[6][18]  = llr_new[6][15];
        llr_in_tmp[6][19]  = llr_new[6][16];
        llr_in_tmp[6][20]  = llr_new[6][17];
        llr_in_tmp[6][21]  = llr_new[6][18];
        llr_in_tmp[6][22]  = llr_new[6][19];
        llr_in_tmp[6][23]  = llr_new[6][20];
        llr_in_tmp[6][24]  = llr_new[6][21];
        llr_in_tmp[6][25]  = llr_new[6][22];
        llr_in_tmp[6][26]  = llr_new[6][23];
        llr_in_tmp[6][27]  = llr_new[6][24];
        llr_in_tmp[6][28]  = llr_new[6][25];
        llr_in_tmp[6][29]  = llr_new[6][26];
        llr_in_tmp[6][30]  = llr_new[6][27];
        llr_in_tmp[6][31]  = llr_new[6][28];
        llr_in_tmp[6][32]  = llr_new[6][29];
        llr_in_tmp[6][33]  = llr_new[6][30];
        llr_in_tmp[6][34]  = llr_new[6][31];
        llr_in_tmp[6][35]  = llr_new[6][32];
        llr_in_tmp[6][36]  = llr_new[6][33];
        llr_in_tmp[6][37]  = llr_new[6][34];
        llr_in_tmp[6][38]  = llr_new[6][35];
        llr_in_tmp[6][39]  = llr_new[6][36];
        llr_in_tmp[6][40]  = llr_new[6][37];
        llr_in_tmp[6][41]  = llr_new[6][38];
    end
 
    5:begin 
        llr_in_tmp[6][0]  = llr_new[6][0];
        llr_in_tmp[6][1]  = llr_new[6][1];
        llr_in_tmp[6][2]  = llr_new[6][2];
        llr_in_tmp[6][3]  = llr_new[6][3];
        llr_in_tmp[6][4]  = llr_new[6][4];
        llr_in_tmp[6][5]  = llr_new[6][5];
        llr_in_tmp[6][6]  = llr_new[6][6];
        llr_in_tmp[6][7]  = llr_new[6][7];
        llr_in_tmp[6][8]  = llr_new[6][8];
        llr_in_tmp[6][9]  = llr_new[6][9];
        llr_in_tmp[6][10]  = llr_new[6][10];
        llr_in_tmp[6][11]  = llr_new[6][11];
        llr_in_tmp[6][12]  = llr_new[6][12];
        llr_in_tmp[6][13]  = llr_new[6][13];
        llr_in_tmp[6][14]  = llr_new[6][14];
        llr_in_tmp[6][15]  = llr_new[6][15];
        llr_in_tmp[6][16]  = llr_new[6][16];
        llr_in_tmp[6][17]  = llr_new[6][17];
        llr_in_tmp[6][18]  = llr_new[6][18];
        llr_in_tmp[6][19]  = llr_new[6][19];
        llr_in_tmp[6][20]  = llr_new[6][20];
        llr_in_tmp[6][21]  = llr_new[6][21];
        llr_in_tmp[6][22]  = llr_new[6][22];
        llr_in_tmp[6][23]  = llr_new[6][23];
        llr_in_tmp[6][24]  = llr_new[6][24];
        llr_in_tmp[6][25]  = llr_new[6][25];
        llr_in_tmp[6][26]  = llr_new[6][26];
        llr_in_tmp[6][27]  = llr_new[6][27];
        llr_in_tmp[6][28]  = llr_new[6][28];
        llr_in_tmp[6][29]  = llr_new[6][29];
        llr_in_tmp[6][30]  = llr_new[6][30];
        llr_in_tmp[6][31]  = llr_new[6][31];
        llr_in_tmp[6][32]  = llr_new[6][32];
        llr_in_tmp[6][33]  = llr_new[6][33];
        llr_in_tmp[6][34]  = llr_new[6][34];
        llr_in_tmp[6][35]  = llr_new[6][35];
        llr_in_tmp[6][36]  = llr_new[6][36];
        llr_in_tmp[6][37]  = llr_new[6][37];
        llr_in_tmp[6][38]  = llr_new[6][38];
        llr_in_tmp[6][39]  = llr_new[6][39];
        llr_in_tmp[6][40]  = llr_new[6][40];
        llr_in_tmp[6][41]  = llr_new[6][41];
    end
 
    6:begin 
        llr_in_tmp[6][0]  = llr_new[6][0];
        llr_in_tmp[6][1]  = llr_new[6][1];
        llr_in_tmp[6][2]  = llr_new[6][2];
        llr_in_tmp[6][3]  = llr_new[6][3];
        llr_in_tmp[6][4]  = llr_new[6][4];
        llr_in_tmp[6][5]  = llr_new[6][5];
        llr_in_tmp[6][6]  = llr_new[6][6];
        llr_in_tmp[6][7]  = llr_new[6][7];
        llr_in_tmp[6][8]  = llr_new[6][8];
        llr_in_tmp[6][9]  = llr_new[6][9];
        llr_in_tmp[6][10]  = llr_new[6][10];
        llr_in_tmp[6][11]  = llr_new[6][11];
        llr_in_tmp[6][12]  = llr_new[6][12];
        llr_in_tmp[6][13]  = llr_new[6][13];
        llr_in_tmp[6][14]  = llr_new[6][14];
        llr_in_tmp[6][15]  = llr_new[6][15];
        llr_in_tmp[6][16]  = llr_new[6][16];
        llr_in_tmp[6][17]  = llr_new[6][17];
        llr_in_tmp[6][18]  = llr_new[6][18];
        llr_in_tmp[6][19]  = llr_new[6][19];
        llr_in_tmp[6][20]  = llr_new[6][20];
        llr_in_tmp[6][21]  = llr_new[6][21];
        llr_in_tmp[6][22]  = llr_new[6][22];
        llr_in_tmp[6][23]  = llr_new[6][23];
        llr_in_tmp[6][24]  = llr_new[6][24];
        llr_in_tmp[6][25]  = llr_new[6][25];
        llr_in_tmp[6][26]  = llr_new[6][26];
        llr_in_tmp[6][27]  = llr_new[6][27];
        llr_in_tmp[6][28]  = llr_new[6][28];
        llr_in_tmp[6][29]  = llr_new[6][29];
        llr_in_tmp[6][30]  = llr_new[6][30];
        llr_in_tmp[6][31]  = llr_new[6][31];
        llr_in_tmp[6][32]  = llr_new[6][32];
        llr_in_tmp[6][33]  = llr_new[6][33];
        llr_in_tmp[6][34]  = llr_new[6][34];
        llr_in_tmp[6][35]  = llr_new[6][35];
        llr_in_tmp[6][36]  = llr_new[6][36];
        llr_in_tmp[6][37]  = llr_new[6][37];
        llr_in_tmp[6][38]  = llr_new[6][38];
        llr_in_tmp[6][39]  = llr_new[6][39];
        llr_in_tmp[6][40]  = llr_new[6][40];
        llr_in_tmp[6][41]  = llr_new[6][41];
    end
 
    7:begin 
        llr_in_tmp[6][0]  = llr_new[6][14];
        llr_in_tmp[6][1]  = llr_new[6][15];
        llr_in_tmp[6][2]  = llr_new[6][16];
        llr_in_tmp[6][3]  = llr_new[6][17];
        llr_in_tmp[6][4]  = llr_new[6][18];
        llr_in_tmp[6][5]  = llr_new[6][19];
        llr_in_tmp[6][6]  = llr_new[6][20];
        llr_in_tmp[6][7]  = llr_new[6][21];
        llr_in_tmp[6][8]  = llr_new[6][22];
        llr_in_tmp[6][9]  = llr_new[6][23];
        llr_in_tmp[6][10]  = llr_new[6][24];
        llr_in_tmp[6][11]  = llr_new[6][25];
        llr_in_tmp[6][12]  = llr_new[6][26];
        llr_in_tmp[6][13]  = llr_new[6][27];
        llr_in_tmp[6][14]  = llr_new[6][28];
        llr_in_tmp[6][15]  = llr_new[6][29];
        llr_in_tmp[6][16]  = llr_new[6][30];
        llr_in_tmp[6][17]  = llr_new[6][31];
        llr_in_tmp[6][18]  = llr_new[6][32];
        llr_in_tmp[6][19]  = llr_new[6][33];
        llr_in_tmp[6][20]  = llr_new[6][34];
        llr_in_tmp[6][21]  = llr_new[6][35];
        llr_in_tmp[6][22]  = llr_new[6][36];
        llr_in_tmp[6][23]  = llr_new[6][37];
        llr_in_tmp[6][24]  = llr_new[6][38];
        llr_in_tmp[6][25]  = llr_new[6][39];
        llr_in_tmp[6][26]  = llr_new[6][40];
        llr_in_tmp[6][27]  = llr_new[6][41];
        llr_in_tmp[6][28]  = llr_new[6][0];
        llr_in_tmp[6][29]  = llr_new[6][1];
        llr_in_tmp[6][30]  = llr_new[6][2];
        llr_in_tmp[6][31]  = llr_new[6][3];
        llr_in_tmp[6][32]  = llr_new[6][4];
        llr_in_tmp[6][33]  = llr_new[6][5];
        llr_in_tmp[6][34]  = llr_new[6][6];
        llr_in_tmp[6][35]  = llr_new[6][7];
        llr_in_tmp[6][36]  = llr_new[6][8];
        llr_in_tmp[6][37]  = llr_new[6][9];
        llr_in_tmp[6][38]  = llr_new[6][10];
        llr_in_tmp[6][39]  = llr_new[6][11];
        llr_in_tmp[6][40]  = llr_new[6][12];
        llr_in_tmp[6][41]  = llr_new[6][13];
    end
 
endcase
end

if (chk_n_input_valid) begin
case (curr_layer)
    0:begin 
        llr_in_tmp[7][0]  = llr_new[7][0];
        llr_in_tmp[7][1]  = llr_new[7][1];
        llr_in_tmp[7][2]  = llr_new[7][2];
        llr_in_tmp[7][3]  = llr_new[7][3];
        llr_in_tmp[7][4]  = llr_new[7][4];
        llr_in_tmp[7][5]  = llr_new[7][5];
        llr_in_tmp[7][6]  = llr_new[7][6];
        llr_in_tmp[7][7]  = llr_new[7][7];
        llr_in_tmp[7][8]  = llr_new[7][8];
        llr_in_tmp[7][9]  = llr_new[7][9];
        llr_in_tmp[7][10]  = llr_new[7][10];
        llr_in_tmp[7][11]  = llr_new[7][11];
        llr_in_tmp[7][12]  = llr_new[7][12];
        llr_in_tmp[7][13]  = llr_new[7][13];
        llr_in_tmp[7][14]  = llr_new[7][14];
        llr_in_tmp[7][15]  = llr_new[7][15];
        llr_in_tmp[7][16]  = llr_new[7][16];
        llr_in_tmp[7][17]  = llr_new[7][17];
        llr_in_tmp[7][18]  = llr_new[7][18];
        llr_in_tmp[7][19]  = llr_new[7][19];
        llr_in_tmp[7][20]  = llr_new[7][20];
        llr_in_tmp[7][21]  = llr_new[7][21];
        llr_in_tmp[7][22]  = llr_new[7][22];
        llr_in_tmp[7][23]  = llr_new[7][23];
        llr_in_tmp[7][24]  = llr_new[7][24];
        llr_in_tmp[7][25]  = llr_new[7][25];
        llr_in_tmp[7][26]  = llr_new[7][26];
        llr_in_tmp[7][27]  = llr_new[7][27];
        llr_in_tmp[7][28]  = llr_new[7][28];
        llr_in_tmp[7][29]  = llr_new[7][29];
        llr_in_tmp[7][30]  = llr_new[7][30];
        llr_in_tmp[7][31]  = llr_new[7][31];
        llr_in_tmp[7][32]  = llr_new[7][32];
        llr_in_tmp[7][33]  = llr_new[7][33];
        llr_in_tmp[7][34]  = llr_new[7][34];
        llr_in_tmp[7][35]  = llr_new[7][35];
        llr_in_tmp[7][36]  = llr_new[7][36];
        llr_in_tmp[7][37]  = llr_new[7][37];
        llr_in_tmp[7][38]  = llr_new[7][38];
        llr_in_tmp[7][39]  = llr_new[7][39];
        llr_in_tmp[7][40]  = llr_new[7][40];
        llr_in_tmp[7][41]  = llr_new[7][41];
    end
 
    1:begin 
        llr_in_tmp[7][0]  = llr_new[7][30];
        llr_in_tmp[7][1]  = llr_new[7][31];
        llr_in_tmp[7][2]  = llr_new[7][32];
        llr_in_tmp[7][3]  = llr_new[7][33];
        llr_in_tmp[7][4]  = llr_new[7][34];
        llr_in_tmp[7][5]  = llr_new[7][35];
        llr_in_tmp[7][6]  = llr_new[7][36];
        llr_in_tmp[7][7]  = llr_new[7][37];
        llr_in_tmp[7][8]  = llr_new[7][38];
        llr_in_tmp[7][9]  = llr_new[7][39];
        llr_in_tmp[7][10]  = llr_new[7][40];
        llr_in_tmp[7][11]  = llr_new[7][41];
        llr_in_tmp[7][12]  = llr_new[7][0];
        llr_in_tmp[7][13]  = llr_new[7][1];
        llr_in_tmp[7][14]  = llr_new[7][2];
        llr_in_tmp[7][15]  = llr_new[7][3];
        llr_in_tmp[7][16]  = llr_new[7][4];
        llr_in_tmp[7][17]  = llr_new[7][5];
        llr_in_tmp[7][18]  = llr_new[7][6];
        llr_in_tmp[7][19]  = llr_new[7][7];
        llr_in_tmp[7][20]  = llr_new[7][8];
        llr_in_tmp[7][21]  = llr_new[7][9];
        llr_in_tmp[7][22]  = llr_new[7][10];
        llr_in_tmp[7][23]  = llr_new[7][11];
        llr_in_tmp[7][24]  = llr_new[7][12];
        llr_in_tmp[7][25]  = llr_new[7][13];
        llr_in_tmp[7][26]  = llr_new[7][14];
        llr_in_tmp[7][27]  = llr_new[7][15];
        llr_in_tmp[7][28]  = llr_new[7][16];
        llr_in_tmp[7][29]  = llr_new[7][17];
        llr_in_tmp[7][30]  = llr_new[7][18];
        llr_in_tmp[7][31]  = llr_new[7][19];
        llr_in_tmp[7][32]  = llr_new[7][20];
        llr_in_tmp[7][33]  = llr_new[7][21];
        llr_in_tmp[7][34]  = llr_new[7][22];
        llr_in_tmp[7][35]  = llr_new[7][23];
        llr_in_tmp[7][36]  = llr_new[7][24];
        llr_in_tmp[7][37]  = llr_new[7][25];
        llr_in_tmp[7][38]  = llr_new[7][26];
        llr_in_tmp[7][39]  = llr_new[7][27];
        llr_in_tmp[7][40]  = llr_new[7][28];
        llr_in_tmp[7][41]  = llr_new[7][29];
    end
 
    2:begin 
        llr_in_tmp[7][0]  = llr_new[7][34];
        llr_in_tmp[7][1]  = llr_new[7][35];
        llr_in_tmp[7][2]  = llr_new[7][36];
        llr_in_tmp[7][3]  = llr_new[7][37];
        llr_in_tmp[7][4]  = llr_new[7][38];
        llr_in_tmp[7][5]  = llr_new[7][39];
        llr_in_tmp[7][6]  = llr_new[7][40];
        llr_in_tmp[7][7]  = llr_new[7][41];
        llr_in_tmp[7][8]  = llr_new[7][0];
        llr_in_tmp[7][9]  = llr_new[7][1];
        llr_in_tmp[7][10]  = llr_new[7][2];
        llr_in_tmp[7][11]  = llr_new[7][3];
        llr_in_tmp[7][12]  = llr_new[7][4];
        llr_in_tmp[7][13]  = llr_new[7][5];
        llr_in_tmp[7][14]  = llr_new[7][6];
        llr_in_tmp[7][15]  = llr_new[7][7];
        llr_in_tmp[7][16]  = llr_new[7][8];
        llr_in_tmp[7][17]  = llr_new[7][9];
        llr_in_tmp[7][18]  = llr_new[7][10];
        llr_in_tmp[7][19]  = llr_new[7][11];
        llr_in_tmp[7][20]  = llr_new[7][12];
        llr_in_tmp[7][21]  = llr_new[7][13];
        llr_in_tmp[7][22]  = llr_new[7][14];
        llr_in_tmp[7][23]  = llr_new[7][15];
        llr_in_tmp[7][24]  = llr_new[7][16];
        llr_in_tmp[7][25]  = llr_new[7][17];
        llr_in_tmp[7][26]  = llr_new[7][18];
        llr_in_tmp[7][27]  = llr_new[7][19];
        llr_in_tmp[7][28]  = llr_new[7][20];
        llr_in_tmp[7][29]  = llr_new[7][21];
        llr_in_tmp[7][30]  = llr_new[7][22];
        llr_in_tmp[7][31]  = llr_new[7][23];
        llr_in_tmp[7][32]  = llr_new[7][24];
        llr_in_tmp[7][33]  = llr_new[7][25];
        llr_in_tmp[7][34]  = llr_new[7][26];
        llr_in_tmp[7][35]  = llr_new[7][27];
        llr_in_tmp[7][36]  = llr_new[7][28];
        llr_in_tmp[7][37]  = llr_new[7][29];
        llr_in_tmp[7][38]  = llr_new[7][30];
        llr_in_tmp[7][39]  = llr_new[7][31];
        llr_in_tmp[7][40]  = llr_new[7][32];
        llr_in_tmp[7][41]  = llr_new[7][33];
    end
 
    3:begin 
        llr_in_tmp[7][0]  = llr_new[7][0];
        llr_in_tmp[7][1]  = llr_new[7][1];
        llr_in_tmp[7][2]  = llr_new[7][2];
        llr_in_tmp[7][3]  = llr_new[7][3];
        llr_in_tmp[7][4]  = llr_new[7][4];
        llr_in_tmp[7][5]  = llr_new[7][5];
        llr_in_tmp[7][6]  = llr_new[7][6];
        llr_in_tmp[7][7]  = llr_new[7][7];
        llr_in_tmp[7][8]  = llr_new[7][8];
        llr_in_tmp[7][9]  = llr_new[7][9];
        llr_in_tmp[7][10]  = llr_new[7][10];
        llr_in_tmp[7][11]  = llr_new[7][11];
        llr_in_tmp[7][12]  = llr_new[7][12];
        llr_in_tmp[7][13]  = llr_new[7][13];
        llr_in_tmp[7][14]  = llr_new[7][14];
        llr_in_tmp[7][15]  = llr_new[7][15];
        llr_in_tmp[7][16]  = llr_new[7][16];
        llr_in_tmp[7][17]  = llr_new[7][17];
        llr_in_tmp[7][18]  = llr_new[7][18];
        llr_in_tmp[7][19]  = llr_new[7][19];
        llr_in_tmp[7][20]  = llr_new[7][20];
        llr_in_tmp[7][21]  = llr_new[7][21];
        llr_in_tmp[7][22]  = llr_new[7][22];
        llr_in_tmp[7][23]  = llr_new[7][23];
        llr_in_tmp[7][24]  = llr_new[7][24];
        llr_in_tmp[7][25]  = llr_new[7][25];
        llr_in_tmp[7][26]  = llr_new[7][26];
        llr_in_tmp[7][27]  = llr_new[7][27];
        llr_in_tmp[7][28]  = llr_new[7][28];
        llr_in_tmp[7][29]  = llr_new[7][29];
        llr_in_tmp[7][30]  = llr_new[7][30];
        llr_in_tmp[7][31]  = llr_new[7][31];
        llr_in_tmp[7][32]  = llr_new[7][32];
        llr_in_tmp[7][33]  = llr_new[7][33];
        llr_in_tmp[7][34]  = llr_new[7][34];
        llr_in_tmp[7][35]  = llr_new[7][35];
        llr_in_tmp[7][36]  = llr_new[7][36];
        llr_in_tmp[7][37]  = llr_new[7][37];
        llr_in_tmp[7][38]  = llr_new[7][38];
        llr_in_tmp[7][39]  = llr_new[7][39];
        llr_in_tmp[7][40]  = llr_new[7][40];
        llr_in_tmp[7][41]  = llr_new[7][41];
    end
 
    4:begin 
        llr_in_tmp[7][0]  = llr_new[7][0];
        llr_in_tmp[7][1]  = llr_new[7][1];
        llr_in_tmp[7][2]  = llr_new[7][2];
        llr_in_tmp[7][3]  = llr_new[7][3];
        llr_in_tmp[7][4]  = llr_new[7][4];
        llr_in_tmp[7][5]  = llr_new[7][5];
        llr_in_tmp[7][6]  = llr_new[7][6];
        llr_in_tmp[7][7]  = llr_new[7][7];
        llr_in_tmp[7][8]  = llr_new[7][8];
        llr_in_tmp[7][9]  = llr_new[7][9];
        llr_in_tmp[7][10]  = llr_new[7][10];
        llr_in_tmp[7][11]  = llr_new[7][11];
        llr_in_tmp[7][12]  = llr_new[7][12];
        llr_in_tmp[7][13]  = llr_new[7][13];
        llr_in_tmp[7][14]  = llr_new[7][14];
        llr_in_tmp[7][15]  = llr_new[7][15];
        llr_in_tmp[7][16]  = llr_new[7][16];
        llr_in_tmp[7][17]  = llr_new[7][17];
        llr_in_tmp[7][18]  = llr_new[7][18];
        llr_in_tmp[7][19]  = llr_new[7][19];
        llr_in_tmp[7][20]  = llr_new[7][20];
        llr_in_tmp[7][21]  = llr_new[7][21];
        llr_in_tmp[7][22]  = llr_new[7][22];
        llr_in_tmp[7][23]  = llr_new[7][23];
        llr_in_tmp[7][24]  = llr_new[7][24];
        llr_in_tmp[7][25]  = llr_new[7][25];
        llr_in_tmp[7][26]  = llr_new[7][26];
        llr_in_tmp[7][27]  = llr_new[7][27];
        llr_in_tmp[7][28]  = llr_new[7][28];
        llr_in_tmp[7][29]  = llr_new[7][29];
        llr_in_tmp[7][30]  = llr_new[7][30];
        llr_in_tmp[7][31]  = llr_new[7][31];
        llr_in_tmp[7][32]  = llr_new[7][32];
        llr_in_tmp[7][33]  = llr_new[7][33];
        llr_in_tmp[7][34]  = llr_new[7][34];
        llr_in_tmp[7][35]  = llr_new[7][35];
        llr_in_tmp[7][36]  = llr_new[7][36];
        llr_in_tmp[7][37]  = llr_new[7][37];
        llr_in_tmp[7][38]  = llr_new[7][38];
        llr_in_tmp[7][39]  = llr_new[7][39];
        llr_in_tmp[7][40]  = llr_new[7][40];
        llr_in_tmp[7][41]  = llr_new[7][41];
    end
 
    5:begin 
        llr_in_tmp[7][0]  = llr_new[7][4];
        llr_in_tmp[7][1]  = llr_new[7][5];
        llr_in_tmp[7][2]  = llr_new[7][6];
        llr_in_tmp[7][3]  = llr_new[7][7];
        llr_in_tmp[7][4]  = llr_new[7][8];
        llr_in_tmp[7][5]  = llr_new[7][9];
        llr_in_tmp[7][6]  = llr_new[7][10];
        llr_in_tmp[7][7]  = llr_new[7][11];
        llr_in_tmp[7][8]  = llr_new[7][12];
        llr_in_tmp[7][9]  = llr_new[7][13];
        llr_in_tmp[7][10]  = llr_new[7][14];
        llr_in_tmp[7][11]  = llr_new[7][15];
        llr_in_tmp[7][12]  = llr_new[7][16];
        llr_in_tmp[7][13]  = llr_new[7][17];
        llr_in_tmp[7][14]  = llr_new[7][18];
        llr_in_tmp[7][15]  = llr_new[7][19];
        llr_in_tmp[7][16]  = llr_new[7][20];
        llr_in_tmp[7][17]  = llr_new[7][21];
        llr_in_tmp[7][18]  = llr_new[7][22];
        llr_in_tmp[7][19]  = llr_new[7][23];
        llr_in_tmp[7][20]  = llr_new[7][24];
        llr_in_tmp[7][21]  = llr_new[7][25];
        llr_in_tmp[7][22]  = llr_new[7][26];
        llr_in_tmp[7][23]  = llr_new[7][27];
        llr_in_tmp[7][24]  = llr_new[7][28];
        llr_in_tmp[7][25]  = llr_new[7][29];
        llr_in_tmp[7][26]  = llr_new[7][30];
        llr_in_tmp[7][27]  = llr_new[7][31];
        llr_in_tmp[7][28]  = llr_new[7][32];
        llr_in_tmp[7][29]  = llr_new[7][33];
        llr_in_tmp[7][30]  = llr_new[7][34];
        llr_in_tmp[7][31]  = llr_new[7][35];
        llr_in_tmp[7][32]  = llr_new[7][36];
        llr_in_tmp[7][33]  = llr_new[7][37];
        llr_in_tmp[7][34]  = llr_new[7][38];
        llr_in_tmp[7][35]  = llr_new[7][39];
        llr_in_tmp[7][36]  = llr_new[7][40];
        llr_in_tmp[7][37]  = llr_new[7][41];
        llr_in_tmp[7][38]  = llr_new[7][0];
        llr_in_tmp[7][39]  = llr_new[7][1];
        llr_in_tmp[7][40]  = llr_new[7][2];
        llr_in_tmp[7][41]  = llr_new[7][3];
    end
 
    6:begin 
        llr_in_tmp[7][0]  = llr_new[7][20];
        llr_in_tmp[7][1]  = llr_new[7][21];
        llr_in_tmp[7][2]  = llr_new[7][22];
        llr_in_tmp[7][3]  = llr_new[7][23];
        llr_in_tmp[7][4]  = llr_new[7][24];
        llr_in_tmp[7][5]  = llr_new[7][25];
        llr_in_tmp[7][6]  = llr_new[7][26];
        llr_in_tmp[7][7]  = llr_new[7][27];
        llr_in_tmp[7][8]  = llr_new[7][28];
        llr_in_tmp[7][9]  = llr_new[7][29];
        llr_in_tmp[7][10]  = llr_new[7][30];
        llr_in_tmp[7][11]  = llr_new[7][31];
        llr_in_tmp[7][12]  = llr_new[7][32];
        llr_in_tmp[7][13]  = llr_new[7][33];
        llr_in_tmp[7][14]  = llr_new[7][34];
        llr_in_tmp[7][15]  = llr_new[7][35];
        llr_in_tmp[7][16]  = llr_new[7][36];
        llr_in_tmp[7][17]  = llr_new[7][37];
        llr_in_tmp[7][18]  = llr_new[7][38];
        llr_in_tmp[7][19]  = llr_new[7][39];
        llr_in_tmp[7][20]  = llr_new[7][40];
        llr_in_tmp[7][21]  = llr_new[7][41];
        llr_in_tmp[7][22]  = llr_new[7][0];
        llr_in_tmp[7][23]  = llr_new[7][1];
        llr_in_tmp[7][24]  = llr_new[7][2];
        llr_in_tmp[7][25]  = llr_new[7][3];
        llr_in_tmp[7][26]  = llr_new[7][4];
        llr_in_tmp[7][27]  = llr_new[7][5];
        llr_in_tmp[7][28]  = llr_new[7][6];
        llr_in_tmp[7][29]  = llr_new[7][7];
        llr_in_tmp[7][30]  = llr_new[7][8];
        llr_in_tmp[7][31]  = llr_new[7][9];
        llr_in_tmp[7][32]  = llr_new[7][10];
        llr_in_tmp[7][33]  = llr_new[7][11];
        llr_in_tmp[7][34]  = llr_new[7][12];
        llr_in_tmp[7][35]  = llr_new[7][13];
        llr_in_tmp[7][36]  = llr_new[7][14];
        llr_in_tmp[7][37]  = llr_new[7][15];
        llr_in_tmp[7][38]  = llr_new[7][16];
        llr_in_tmp[7][39]  = llr_new[7][17];
        llr_in_tmp[7][40]  = llr_new[7][18];
        llr_in_tmp[7][41]  = llr_new[7][19];
    end
 
    7:begin 
        llr_in_tmp[7][0]  = llr_new[7][0];
        llr_in_tmp[7][1]  = llr_new[7][1];
        llr_in_tmp[7][2]  = llr_new[7][2];
        llr_in_tmp[7][3]  = llr_new[7][3];
        llr_in_tmp[7][4]  = llr_new[7][4];
        llr_in_tmp[7][5]  = llr_new[7][5];
        llr_in_tmp[7][6]  = llr_new[7][6];
        llr_in_tmp[7][7]  = llr_new[7][7];
        llr_in_tmp[7][8]  = llr_new[7][8];
        llr_in_tmp[7][9]  = llr_new[7][9];
        llr_in_tmp[7][10]  = llr_new[7][10];
        llr_in_tmp[7][11]  = llr_new[7][11];
        llr_in_tmp[7][12]  = llr_new[7][12];
        llr_in_tmp[7][13]  = llr_new[7][13];
        llr_in_tmp[7][14]  = llr_new[7][14];
        llr_in_tmp[7][15]  = llr_new[7][15];
        llr_in_tmp[7][16]  = llr_new[7][16];
        llr_in_tmp[7][17]  = llr_new[7][17];
        llr_in_tmp[7][18]  = llr_new[7][18];
        llr_in_tmp[7][19]  = llr_new[7][19];
        llr_in_tmp[7][20]  = llr_new[7][20];
        llr_in_tmp[7][21]  = llr_new[7][21];
        llr_in_tmp[7][22]  = llr_new[7][22];
        llr_in_tmp[7][23]  = llr_new[7][23];
        llr_in_tmp[7][24]  = llr_new[7][24];
        llr_in_tmp[7][25]  = llr_new[7][25];
        llr_in_tmp[7][26]  = llr_new[7][26];
        llr_in_tmp[7][27]  = llr_new[7][27];
        llr_in_tmp[7][28]  = llr_new[7][28];
        llr_in_tmp[7][29]  = llr_new[7][29];
        llr_in_tmp[7][30]  = llr_new[7][30];
        llr_in_tmp[7][31]  = llr_new[7][31];
        llr_in_tmp[7][32]  = llr_new[7][32];
        llr_in_tmp[7][33]  = llr_new[7][33];
        llr_in_tmp[7][34]  = llr_new[7][34];
        llr_in_tmp[7][35]  = llr_new[7][35];
        llr_in_tmp[7][36]  = llr_new[7][36];
        llr_in_tmp[7][37]  = llr_new[7][37];
        llr_in_tmp[7][38]  = llr_new[7][38];
        llr_in_tmp[7][39]  = llr_new[7][39];
        llr_in_tmp[7][40]  = llr_new[7][40];
        llr_in_tmp[7][41]  = llr_new[7][41];
    end
 
endcase
end

if (chk_n_input_valid) begin
case (curr_layer)
    0:begin 
        llr_in_tmp[8][0]  = llr_new[8][18];
        llr_in_tmp[8][1]  = llr_new[8][19];
        llr_in_tmp[8][2]  = llr_new[8][20];
        llr_in_tmp[8][3]  = llr_new[8][21];
        llr_in_tmp[8][4]  = llr_new[8][22];
        llr_in_tmp[8][5]  = llr_new[8][23];
        llr_in_tmp[8][6]  = llr_new[8][24];
        llr_in_tmp[8][7]  = llr_new[8][25];
        llr_in_tmp[8][8]  = llr_new[8][26];
        llr_in_tmp[8][9]  = llr_new[8][27];
        llr_in_tmp[8][10]  = llr_new[8][28];
        llr_in_tmp[8][11]  = llr_new[8][29];
        llr_in_tmp[8][12]  = llr_new[8][30];
        llr_in_tmp[8][13]  = llr_new[8][31];
        llr_in_tmp[8][14]  = llr_new[8][32];
        llr_in_tmp[8][15]  = llr_new[8][33];
        llr_in_tmp[8][16]  = llr_new[8][34];
        llr_in_tmp[8][17]  = llr_new[8][35];
        llr_in_tmp[8][18]  = llr_new[8][36];
        llr_in_tmp[8][19]  = llr_new[8][37];
        llr_in_tmp[8][20]  = llr_new[8][38];
        llr_in_tmp[8][21]  = llr_new[8][39];
        llr_in_tmp[8][22]  = llr_new[8][40];
        llr_in_tmp[8][23]  = llr_new[8][41];
        llr_in_tmp[8][24]  = llr_new[8][0];
        llr_in_tmp[8][25]  = llr_new[8][1];
        llr_in_tmp[8][26]  = llr_new[8][2];
        llr_in_tmp[8][27]  = llr_new[8][3];
        llr_in_tmp[8][28]  = llr_new[8][4];
        llr_in_tmp[8][29]  = llr_new[8][5];
        llr_in_tmp[8][30]  = llr_new[8][6];
        llr_in_tmp[8][31]  = llr_new[8][7];
        llr_in_tmp[8][32]  = llr_new[8][8];
        llr_in_tmp[8][33]  = llr_new[8][9];
        llr_in_tmp[8][34]  = llr_new[8][10];
        llr_in_tmp[8][35]  = llr_new[8][11];
        llr_in_tmp[8][36]  = llr_new[8][12];
        llr_in_tmp[8][37]  = llr_new[8][13];
        llr_in_tmp[8][38]  = llr_new[8][14];
        llr_in_tmp[8][39]  = llr_new[8][15];
        llr_in_tmp[8][40]  = llr_new[8][16];
        llr_in_tmp[8][41]  = llr_new[8][17];
    end
 
    1:begin 
        llr_in_tmp[8][0]  = llr_new[8][2];
        llr_in_tmp[8][1]  = llr_new[8][3];
        llr_in_tmp[8][2]  = llr_new[8][4];
        llr_in_tmp[8][3]  = llr_new[8][5];
        llr_in_tmp[8][4]  = llr_new[8][6];
        llr_in_tmp[8][5]  = llr_new[8][7];
        llr_in_tmp[8][6]  = llr_new[8][8];
        llr_in_tmp[8][7]  = llr_new[8][9];
        llr_in_tmp[8][8]  = llr_new[8][10];
        llr_in_tmp[8][9]  = llr_new[8][11];
        llr_in_tmp[8][10]  = llr_new[8][12];
        llr_in_tmp[8][11]  = llr_new[8][13];
        llr_in_tmp[8][12]  = llr_new[8][14];
        llr_in_tmp[8][13]  = llr_new[8][15];
        llr_in_tmp[8][14]  = llr_new[8][16];
        llr_in_tmp[8][15]  = llr_new[8][17];
        llr_in_tmp[8][16]  = llr_new[8][18];
        llr_in_tmp[8][17]  = llr_new[8][19];
        llr_in_tmp[8][18]  = llr_new[8][20];
        llr_in_tmp[8][19]  = llr_new[8][21];
        llr_in_tmp[8][20]  = llr_new[8][22];
        llr_in_tmp[8][21]  = llr_new[8][23];
        llr_in_tmp[8][22]  = llr_new[8][24];
        llr_in_tmp[8][23]  = llr_new[8][25];
        llr_in_tmp[8][24]  = llr_new[8][26];
        llr_in_tmp[8][25]  = llr_new[8][27];
        llr_in_tmp[8][26]  = llr_new[8][28];
        llr_in_tmp[8][27]  = llr_new[8][29];
        llr_in_tmp[8][28]  = llr_new[8][30];
        llr_in_tmp[8][29]  = llr_new[8][31];
        llr_in_tmp[8][30]  = llr_new[8][32];
        llr_in_tmp[8][31]  = llr_new[8][33];
        llr_in_tmp[8][32]  = llr_new[8][34];
        llr_in_tmp[8][33]  = llr_new[8][35];
        llr_in_tmp[8][34]  = llr_new[8][36];
        llr_in_tmp[8][35]  = llr_new[8][37];
        llr_in_tmp[8][36]  = llr_new[8][38];
        llr_in_tmp[8][37]  = llr_new[8][39];
        llr_in_tmp[8][38]  = llr_new[8][40];
        llr_in_tmp[8][39]  = llr_new[8][41];
        llr_in_tmp[8][40]  = llr_new[8][0];
        llr_in_tmp[8][41]  = llr_new[8][1];
    end
 
    2:begin 
        llr_in_tmp[8][0]  = llr_new[8][0];
        llr_in_tmp[8][1]  = llr_new[8][1];
        llr_in_tmp[8][2]  = llr_new[8][2];
        llr_in_tmp[8][3]  = llr_new[8][3];
        llr_in_tmp[8][4]  = llr_new[8][4];
        llr_in_tmp[8][5]  = llr_new[8][5];
        llr_in_tmp[8][6]  = llr_new[8][6];
        llr_in_tmp[8][7]  = llr_new[8][7];
        llr_in_tmp[8][8]  = llr_new[8][8];
        llr_in_tmp[8][9]  = llr_new[8][9];
        llr_in_tmp[8][10]  = llr_new[8][10];
        llr_in_tmp[8][11]  = llr_new[8][11];
        llr_in_tmp[8][12]  = llr_new[8][12];
        llr_in_tmp[8][13]  = llr_new[8][13];
        llr_in_tmp[8][14]  = llr_new[8][14];
        llr_in_tmp[8][15]  = llr_new[8][15];
        llr_in_tmp[8][16]  = llr_new[8][16];
        llr_in_tmp[8][17]  = llr_new[8][17];
        llr_in_tmp[8][18]  = llr_new[8][18];
        llr_in_tmp[8][19]  = llr_new[8][19];
        llr_in_tmp[8][20]  = llr_new[8][20];
        llr_in_tmp[8][21]  = llr_new[8][21];
        llr_in_tmp[8][22]  = llr_new[8][22];
        llr_in_tmp[8][23]  = llr_new[8][23];
        llr_in_tmp[8][24]  = llr_new[8][24];
        llr_in_tmp[8][25]  = llr_new[8][25];
        llr_in_tmp[8][26]  = llr_new[8][26];
        llr_in_tmp[8][27]  = llr_new[8][27];
        llr_in_tmp[8][28]  = llr_new[8][28];
        llr_in_tmp[8][29]  = llr_new[8][29];
        llr_in_tmp[8][30]  = llr_new[8][30];
        llr_in_tmp[8][31]  = llr_new[8][31];
        llr_in_tmp[8][32]  = llr_new[8][32];
        llr_in_tmp[8][33]  = llr_new[8][33];
        llr_in_tmp[8][34]  = llr_new[8][34];
        llr_in_tmp[8][35]  = llr_new[8][35];
        llr_in_tmp[8][36]  = llr_new[8][36];
        llr_in_tmp[8][37]  = llr_new[8][37];
        llr_in_tmp[8][38]  = llr_new[8][38];
        llr_in_tmp[8][39]  = llr_new[8][39];
        llr_in_tmp[8][40]  = llr_new[8][40];
        llr_in_tmp[8][41]  = llr_new[8][41];
    end
 
    3:begin 
        llr_in_tmp[8][0]  = llr_new[8][0];
        llr_in_tmp[8][1]  = llr_new[8][1];
        llr_in_tmp[8][2]  = llr_new[8][2];
        llr_in_tmp[8][3]  = llr_new[8][3];
        llr_in_tmp[8][4]  = llr_new[8][4];
        llr_in_tmp[8][5]  = llr_new[8][5];
        llr_in_tmp[8][6]  = llr_new[8][6];
        llr_in_tmp[8][7]  = llr_new[8][7];
        llr_in_tmp[8][8]  = llr_new[8][8];
        llr_in_tmp[8][9]  = llr_new[8][9];
        llr_in_tmp[8][10]  = llr_new[8][10];
        llr_in_tmp[8][11]  = llr_new[8][11];
        llr_in_tmp[8][12]  = llr_new[8][12];
        llr_in_tmp[8][13]  = llr_new[8][13];
        llr_in_tmp[8][14]  = llr_new[8][14];
        llr_in_tmp[8][15]  = llr_new[8][15];
        llr_in_tmp[8][16]  = llr_new[8][16];
        llr_in_tmp[8][17]  = llr_new[8][17];
        llr_in_tmp[8][18]  = llr_new[8][18];
        llr_in_tmp[8][19]  = llr_new[8][19];
        llr_in_tmp[8][20]  = llr_new[8][20];
        llr_in_tmp[8][21]  = llr_new[8][21];
        llr_in_tmp[8][22]  = llr_new[8][22];
        llr_in_tmp[8][23]  = llr_new[8][23];
        llr_in_tmp[8][24]  = llr_new[8][24];
        llr_in_tmp[8][25]  = llr_new[8][25];
        llr_in_tmp[8][26]  = llr_new[8][26];
        llr_in_tmp[8][27]  = llr_new[8][27];
        llr_in_tmp[8][28]  = llr_new[8][28];
        llr_in_tmp[8][29]  = llr_new[8][29];
        llr_in_tmp[8][30]  = llr_new[8][30];
        llr_in_tmp[8][31]  = llr_new[8][31];
        llr_in_tmp[8][32]  = llr_new[8][32];
        llr_in_tmp[8][33]  = llr_new[8][33];
        llr_in_tmp[8][34]  = llr_new[8][34];
        llr_in_tmp[8][35]  = llr_new[8][35];
        llr_in_tmp[8][36]  = llr_new[8][36];
        llr_in_tmp[8][37]  = llr_new[8][37];
        llr_in_tmp[8][38]  = llr_new[8][38];
        llr_in_tmp[8][39]  = llr_new[8][39];
        llr_in_tmp[8][40]  = llr_new[8][40];
        llr_in_tmp[8][41]  = llr_new[8][41];
    end
 
    4:begin 
        llr_in_tmp[8][0]  = llr_new[8][28];
        llr_in_tmp[8][1]  = llr_new[8][29];
        llr_in_tmp[8][2]  = llr_new[8][30];
        llr_in_tmp[8][3]  = llr_new[8][31];
        llr_in_tmp[8][4]  = llr_new[8][32];
        llr_in_tmp[8][5]  = llr_new[8][33];
        llr_in_tmp[8][6]  = llr_new[8][34];
        llr_in_tmp[8][7]  = llr_new[8][35];
        llr_in_tmp[8][8]  = llr_new[8][36];
        llr_in_tmp[8][9]  = llr_new[8][37];
        llr_in_tmp[8][10]  = llr_new[8][38];
        llr_in_tmp[8][11]  = llr_new[8][39];
        llr_in_tmp[8][12]  = llr_new[8][40];
        llr_in_tmp[8][13]  = llr_new[8][41];
        llr_in_tmp[8][14]  = llr_new[8][0];
        llr_in_tmp[8][15]  = llr_new[8][1];
        llr_in_tmp[8][16]  = llr_new[8][2];
        llr_in_tmp[8][17]  = llr_new[8][3];
        llr_in_tmp[8][18]  = llr_new[8][4];
        llr_in_tmp[8][19]  = llr_new[8][5];
        llr_in_tmp[8][20]  = llr_new[8][6];
        llr_in_tmp[8][21]  = llr_new[8][7];
        llr_in_tmp[8][22]  = llr_new[8][8];
        llr_in_tmp[8][23]  = llr_new[8][9];
        llr_in_tmp[8][24]  = llr_new[8][10];
        llr_in_tmp[8][25]  = llr_new[8][11];
        llr_in_tmp[8][26]  = llr_new[8][12];
        llr_in_tmp[8][27]  = llr_new[8][13];
        llr_in_tmp[8][28]  = llr_new[8][14];
        llr_in_tmp[8][29]  = llr_new[8][15];
        llr_in_tmp[8][30]  = llr_new[8][16];
        llr_in_tmp[8][31]  = llr_new[8][17];
        llr_in_tmp[8][32]  = llr_new[8][18];
        llr_in_tmp[8][33]  = llr_new[8][19];
        llr_in_tmp[8][34]  = llr_new[8][20];
        llr_in_tmp[8][35]  = llr_new[8][21];
        llr_in_tmp[8][36]  = llr_new[8][22];
        llr_in_tmp[8][37]  = llr_new[8][23];
        llr_in_tmp[8][38]  = llr_new[8][24];
        llr_in_tmp[8][39]  = llr_new[8][25];
        llr_in_tmp[8][40]  = llr_new[8][26];
        llr_in_tmp[8][41]  = llr_new[8][27];
    end
 
    5:begin 
        llr_in_tmp[8][0]  = llr_new[8][0];
        llr_in_tmp[8][1]  = llr_new[8][1];
        llr_in_tmp[8][2]  = llr_new[8][2];
        llr_in_tmp[8][3]  = llr_new[8][3];
        llr_in_tmp[8][4]  = llr_new[8][4];
        llr_in_tmp[8][5]  = llr_new[8][5];
        llr_in_tmp[8][6]  = llr_new[8][6];
        llr_in_tmp[8][7]  = llr_new[8][7];
        llr_in_tmp[8][8]  = llr_new[8][8];
        llr_in_tmp[8][9]  = llr_new[8][9];
        llr_in_tmp[8][10]  = llr_new[8][10];
        llr_in_tmp[8][11]  = llr_new[8][11];
        llr_in_tmp[8][12]  = llr_new[8][12];
        llr_in_tmp[8][13]  = llr_new[8][13];
        llr_in_tmp[8][14]  = llr_new[8][14];
        llr_in_tmp[8][15]  = llr_new[8][15];
        llr_in_tmp[8][16]  = llr_new[8][16];
        llr_in_tmp[8][17]  = llr_new[8][17];
        llr_in_tmp[8][18]  = llr_new[8][18];
        llr_in_tmp[8][19]  = llr_new[8][19];
        llr_in_tmp[8][20]  = llr_new[8][20];
        llr_in_tmp[8][21]  = llr_new[8][21];
        llr_in_tmp[8][22]  = llr_new[8][22];
        llr_in_tmp[8][23]  = llr_new[8][23];
        llr_in_tmp[8][24]  = llr_new[8][24];
        llr_in_tmp[8][25]  = llr_new[8][25];
        llr_in_tmp[8][26]  = llr_new[8][26];
        llr_in_tmp[8][27]  = llr_new[8][27];
        llr_in_tmp[8][28]  = llr_new[8][28];
        llr_in_tmp[8][29]  = llr_new[8][29];
        llr_in_tmp[8][30]  = llr_new[8][30];
        llr_in_tmp[8][31]  = llr_new[8][31];
        llr_in_tmp[8][32]  = llr_new[8][32];
        llr_in_tmp[8][33]  = llr_new[8][33];
        llr_in_tmp[8][34]  = llr_new[8][34];
        llr_in_tmp[8][35]  = llr_new[8][35];
        llr_in_tmp[8][36]  = llr_new[8][36];
        llr_in_tmp[8][37]  = llr_new[8][37];
        llr_in_tmp[8][38]  = llr_new[8][38];
        llr_in_tmp[8][39]  = llr_new[8][39];
        llr_in_tmp[8][40]  = llr_new[8][40];
        llr_in_tmp[8][41]  = llr_new[8][41];
    end
 
    6:begin 
        llr_in_tmp[8][0]  = llr_new[8][0];
        llr_in_tmp[8][1]  = llr_new[8][1];
        llr_in_tmp[8][2]  = llr_new[8][2];
        llr_in_tmp[8][3]  = llr_new[8][3];
        llr_in_tmp[8][4]  = llr_new[8][4];
        llr_in_tmp[8][5]  = llr_new[8][5];
        llr_in_tmp[8][6]  = llr_new[8][6];
        llr_in_tmp[8][7]  = llr_new[8][7];
        llr_in_tmp[8][8]  = llr_new[8][8];
        llr_in_tmp[8][9]  = llr_new[8][9];
        llr_in_tmp[8][10]  = llr_new[8][10];
        llr_in_tmp[8][11]  = llr_new[8][11];
        llr_in_tmp[8][12]  = llr_new[8][12];
        llr_in_tmp[8][13]  = llr_new[8][13];
        llr_in_tmp[8][14]  = llr_new[8][14];
        llr_in_tmp[8][15]  = llr_new[8][15];
        llr_in_tmp[8][16]  = llr_new[8][16];
        llr_in_tmp[8][17]  = llr_new[8][17];
        llr_in_tmp[8][18]  = llr_new[8][18];
        llr_in_tmp[8][19]  = llr_new[8][19];
        llr_in_tmp[8][20]  = llr_new[8][20];
        llr_in_tmp[8][21]  = llr_new[8][21];
        llr_in_tmp[8][22]  = llr_new[8][22];
        llr_in_tmp[8][23]  = llr_new[8][23];
        llr_in_tmp[8][24]  = llr_new[8][24];
        llr_in_tmp[8][25]  = llr_new[8][25];
        llr_in_tmp[8][26]  = llr_new[8][26];
        llr_in_tmp[8][27]  = llr_new[8][27];
        llr_in_tmp[8][28]  = llr_new[8][28];
        llr_in_tmp[8][29]  = llr_new[8][29];
        llr_in_tmp[8][30]  = llr_new[8][30];
        llr_in_tmp[8][31]  = llr_new[8][31];
        llr_in_tmp[8][32]  = llr_new[8][32];
        llr_in_tmp[8][33]  = llr_new[8][33];
        llr_in_tmp[8][34]  = llr_new[8][34];
        llr_in_tmp[8][35]  = llr_new[8][35];
        llr_in_tmp[8][36]  = llr_new[8][36];
        llr_in_tmp[8][37]  = llr_new[8][37];
        llr_in_tmp[8][38]  = llr_new[8][38];
        llr_in_tmp[8][39]  = llr_new[8][39];
        llr_in_tmp[8][40]  = llr_new[8][40];
        llr_in_tmp[8][41]  = llr_new[8][41];
    end
 
    7:begin 
        llr_in_tmp[8][0]  = llr_new[8][4];
        llr_in_tmp[8][1]  = llr_new[8][5];
        llr_in_tmp[8][2]  = llr_new[8][6];
        llr_in_tmp[8][3]  = llr_new[8][7];
        llr_in_tmp[8][4]  = llr_new[8][8];
        llr_in_tmp[8][5]  = llr_new[8][9];
        llr_in_tmp[8][6]  = llr_new[8][10];
        llr_in_tmp[8][7]  = llr_new[8][11];
        llr_in_tmp[8][8]  = llr_new[8][12];
        llr_in_tmp[8][9]  = llr_new[8][13];
        llr_in_tmp[8][10]  = llr_new[8][14];
        llr_in_tmp[8][11]  = llr_new[8][15];
        llr_in_tmp[8][12]  = llr_new[8][16];
        llr_in_tmp[8][13]  = llr_new[8][17];
        llr_in_tmp[8][14]  = llr_new[8][18];
        llr_in_tmp[8][15]  = llr_new[8][19];
        llr_in_tmp[8][16]  = llr_new[8][20];
        llr_in_tmp[8][17]  = llr_new[8][21];
        llr_in_tmp[8][18]  = llr_new[8][22];
        llr_in_tmp[8][19]  = llr_new[8][23];
        llr_in_tmp[8][20]  = llr_new[8][24];
        llr_in_tmp[8][21]  = llr_new[8][25];
        llr_in_tmp[8][22]  = llr_new[8][26];
        llr_in_tmp[8][23]  = llr_new[8][27];
        llr_in_tmp[8][24]  = llr_new[8][28];
        llr_in_tmp[8][25]  = llr_new[8][29];
        llr_in_tmp[8][26]  = llr_new[8][30];
        llr_in_tmp[8][27]  = llr_new[8][31];
        llr_in_tmp[8][28]  = llr_new[8][32];
        llr_in_tmp[8][29]  = llr_new[8][33];
        llr_in_tmp[8][30]  = llr_new[8][34];
        llr_in_tmp[8][31]  = llr_new[8][35];
        llr_in_tmp[8][32]  = llr_new[8][36];
        llr_in_tmp[8][33]  = llr_new[8][37];
        llr_in_tmp[8][34]  = llr_new[8][38];
        llr_in_tmp[8][35]  = llr_new[8][39];
        llr_in_tmp[8][36]  = llr_new[8][40];
        llr_in_tmp[8][37]  = llr_new[8][41];
        llr_in_tmp[8][38]  = llr_new[8][0];
        llr_in_tmp[8][39]  = llr_new[8][1];
        llr_in_tmp[8][40]  = llr_new[8][2];
        llr_in_tmp[8][41]  = llr_new[8][3];
    end
 
endcase
end

if (chk_n_input_valid) begin
case (curr_layer)
    0:begin 
        llr_in_tmp[9][0]  = llr_new[9][0];
        llr_in_tmp[9][1]  = llr_new[9][1];
        llr_in_tmp[9][2]  = llr_new[9][2];
        llr_in_tmp[9][3]  = llr_new[9][3];
        llr_in_tmp[9][4]  = llr_new[9][4];
        llr_in_tmp[9][5]  = llr_new[9][5];
        llr_in_tmp[9][6]  = llr_new[9][6];
        llr_in_tmp[9][7]  = llr_new[9][7];
        llr_in_tmp[9][8]  = llr_new[9][8];
        llr_in_tmp[9][9]  = llr_new[9][9];
        llr_in_tmp[9][10]  = llr_new[9][10];
        llr_in_tmp[9][11]  = llr_new[9][11];
        llr_in_tmp[9][12]  = llr_new[9][12];
        llr_in_tmp[9][13]  = llr_new[9][13];
        llr_in_tmp[9][14]  = llr_new[9][14];
        llr_in_tmp[9][15]  = llr_new[9][15];
        llr_in_tmp[9][16]  = llr_new[9][16];
        llr_in_tmp[9][17]  = llr_new[9][17];
        llr_in_tmp[9][18]  = llr_new[9][18];
        llr_in_tmp[9][19]  = llr_new[9][19];
        llr_in_tmp[9][20]  = llr_new[9][20];
        llr_in_tmp[9][21]  = llr_new[9][21];
        llr_in_tmp[9][22]  = llr_new[9][22];
        llr_in_tmp[9][23]  = llr_new[9][23];
        llr_in_tmp[9][24]  = llr_new[9][24];
        llr_in_tmp[9][25]  = llr_new[9][25];
        llr_in_tmp[9][26]  = llr_new[9][26];
        llr_in_tmp[9][27]  = llr_new[9][27];
        llr_in_tmp[9][28]  = llr_new[9][28];
        llr_in_tmp[9][29]  = llr_new[9][29];
        llr_in_tmp[9][30]  = llr_new[9][30];
        llr_in_tmp[9][31]  = llr_new[9][31];
        llr_in_tmp[9][32]  = llr_new[9][32];
        llr_in_tmp[9][33]  = llr_new[9][33];
        llr_in_tmp[9][34]  = llr_new[9][34];
        llr_in_tmp[9][35]  = llr_new[9][35];
        llr_in_tmp[9][36]  = llr_new[9][36];
        llr_in_tmp[9][37]  = llr_new[9][37];
        llr_in_tmp[9][38]  = llr_new[9][38];
        llr_in_tmp[9][39]  = llr_new[9][39];
        llr_in_tmp[9][40]  = llr_new[9][40];
        llr_in_tmp[9][41]  = llr_new[9][41];
    end
 
    1:begin 
        llr_in_tmp[9][0]  = llr_new[9][1];
        llr_in_tmp[9][1]  = llr_new[9][2];
        llr_in_tmp[9][2]  = llr_new[9][3];
        llr_in_tmp[9][3]  = llr_new[9][4];
        llr_in_tmp[9][4]  = llr_new[9][5];
        llr_in_tmp[9][5]  = llr_new[9][6];
        llr_in_tmp[9][6]  = llr_new[9][7];
        llr_in_tmp[9][7]  = llr_new[9][8];
        llr_in_tmp[9][8]  = llr_new[9][9];
        llr_in_tmp[9][9]  = llr_new[9][10];
        llr_in_tmp[9][10]  = llr_new[9][11];
        llr_in_tmp[9][11]  = llr_new[9][12];
        llr_in_tmp[9][12]  = llr_new[9][13];
        llr_in_tmp[9][13]  = llr_new[9][14];
        llr_in_tmp[9][14]  = llr_new[9][15];
        llr_in_tmp[9][15]  = llr_new[9][16];
        llr_in_tmp[9][16]  = llr_new[9][17];
        llr_in_tmp[9][17]  = llr_new[9][18];
        llr_in_tmp[9][18]  = llr_new[9][19];
        llr_in_tmp[9][19]  = llr_new[9][20];
        llr_in_tmp[9][20]  = llr_new[9][21];
        llr_in_tmp[9][21]  = llr_new[9][22];
        llr_in_tmp[9][22]  = llr_new[9][23];
        llr_in_tmp[9][23]  = llr_new[9][24];
        llr_in_tmp[9][24]  = llr_new[9][25];
        llr_in_tmp[9][25]  = llr_new[9][26];
        llr_in_tmp[9][26]  = llr_new[9][27];
        llr_in_tmp[9][27]  = llr_new[9][28];
        llr_in_tmp[9][28]  = llr_new[9][29];
        llr_in_tmp[9][29]  = llr_new[9][30];
        llr_in_tmp[9][30]  = llr_new[9][31];
        llr_in_tmp[9][31]  = llr_new[9][32];
        llr_in_tmp[9][32]  = llr_new[9][33];
        llr_in_tmp[9][33]  = llr_new[9][34];
        llr_in_tmp[9][34]  = llr_new[9][35];
        llr_in_tmp[9][35]  = llr_new[9][36];
        llr_in_tmp[9][36]  = llr_new[9][37];
        llr_in_tmp[9][37]  = llr_new[9][38];
        llr_in_tmp[9][38]  = llr_new[9][39];
        llr_in_tmp[9][39]  = llr_new[9][40];
        llr_in_tmp[9][40]  = llr_new[9][41];
        llr_in_tmp[9][41]  = llr_new[9][0];
    end
 
    2:begin 
        llr_in_tmp[9][0]  = llr_new[9][10];
        llr_in_tmp[9][1]  = llr_new[9][11];
        llr_in_tmp[9][2]  = llr_new[9][12];
        llr_in_tmp[9][3]  = llr_new[9][13];
        llr_in_tmp[9][4]  = llr_new[9][14];
        llr_in_tmp[9][5]  = llr_new[9][15];
        llr_in_tmp[9][6]  = llr_new[9][16];
        llr_in_tmp[9][7]  = llr_new[9][17];
        llr_in_tmp[9][8]  = llr_new[9][18];
        llr_in_tmp[9][9]  = llr_new[9][19];
        llr_in_tmp[9][10]  = llr_new[9][20];
        llr_in_tmp[9][11]  = llr_new[9][21];
        llr_in_tmp[9][12]  = llr_new[9][22];
        llr_in_tmp[9][13]  = llr_new[9][23];
        llr_in_tmp[9][14]  = llr_new[9][24];
        llr_in_tmp[9][15]  = llr_new[9][25];
        llr_in_tmp[9][16]  = llr_new[9][26];
        llr_in_tmp[9][17]  = llr_new[9][27];
        llr_in_tmp[9][18]  = llr_new[9][28];
        llr_in_tmp[9][19]  = llr_new[9][29];
        llr_in_tmp[9][20]  = llr_new[9][30];
        llr_in_tmp[9][21]  = llr_new[9][31];
        llr_in_tmp[9][22]  = llr_new[9][32];
        llr_in_tmp[9][23]  = llr_new[9][33];
        llr_in_tmp[9][24]  = llr_new[9][34];
        llr_in_tmp[9][25]  = llr_new[9][35];
        llr_in_tmp[9][26]  = llr_new[9][36];
        llr_in_tmp[9][27]  = llr_new[9][37];
        llr_in_tmp[9][28]  = llr_new[9][38];
        llr_in_tmp[9][29]  = llr_new[9][39];
        llr_in_tmp[9][30]  = llr_new[9][40];
        llr_in_tmp[9][31]  = llr_new[9][41];
        llr_in_tmp[9][32]  = llr_new[9][0];
        llr_in_tmp[9][33]  = llr_new[9][1];
        llr_in_tmp[9][34]  = llr_new[9][2];
        llr_in_tmp[9][35]  = llr_new[9][3];
        llr_in_tmp[9][36]  = llr_new[9][4];
        llr_in_tmp[9][37]  = llr_new[9][5];
        llr_in_tmp[9][38]  = llr_new[9][6];
        llr_in_tmp[9][39]  = llr_new[9][7];
        llr_in_tmp[9][40]  = llr_new[9][8];
        llr_in_tmp[9][41]  = llr_new[9][9];
    end
 
    3:begin 
        llr_in_tmp[9][0]  = llr_new[9][0];
        llr_in_tmp[9][1]  = llr_new[9][1];
        llr_in_tmp[9][2]  = llr_new[9][2];
        llr_in_tmp[9][3]  = llr_new[9][3];
        llr_in_tmp[9][4]  = llr_new[9][4];
        llr_in_tmp[9][5]  = llr_new[9][5];
        llr_in_tmp[9][6]  = llr_new[9][6];
        llr_in_tmp[9][7]  = llr_new[9][7];
        llr_in_tmp[9][8]  = llr_new[9][8];
        llr_in_tmp[9][9]  = llr_new[9][9];
        llr_in_tmp[9][10]  = llr_new[9][10];
        llr_in_tmp[9][11]  = llr_new[9][11];
        llr_in_tmp[9][12]  = llr_new[9][12];
        llr_in_tmp[9][13]  = llr_new[9][13];
        llr_in_tmp[9][14]  = llr_new[9][14];
        llr_in_tmp[9][15]  = llr_new[9][15];
        llr_in_tmp[9][16]  = llr_new[9][16];
        llr_in_tmp[9][17]  = llr_new[9][17];
        llr_in_tmp[9][18]  = llr_new[9][18];
        llr_in_tmp[9][19]  = llr_new[9][19];
        llr_in_tmp[9][20]  = llr_new[9][20];
        llr_in_tmp[9][21]  = llr_new[9][21];
        llr_in_tmp[9][22]  = llr_new[9][22];
        llr_in_tmp[9][23]  = llr_new[9][23];
        llr_in_tmp[9][24]  = llr_new[9][24];
        llr_in_tmp[9][25]  = llr_new[9][25];
        llr_in_tmp[9][26]  = llr_new[9][26];
        llr_in_tmp[9][27]  = llr_new[9][27];
        llr_in_tmp[9][28]  = llr_new[9][28];
        llr_in_tmp[9][29]  = llr_new[9][29];
        llr_in_tmp[9][30]  = llr_new[9][30];
        llr_in_tmp[9][31]  = llr_new[9][31];
        llr_in_tmp[9][32]  = llr_new[9][32];
        llr_in_tmp[9][33]  = llr_new[9][33];
        llr_in_tmp[9][34]  = llr_new[9][34];
        llr_in_tmp[9][35]  = llr_new[9][35];
        llr_in_tmp[9][36]  = llr_new[9][36];
        llr_in_tmp[9][37]  = llr_new[9][37];
        llr_in_tmp[9][38]  = llr_new[9][38];
        llr_in_tmp[9][39]  = llr_new[9][39];
        llr_in_tmp[9][40]  = llr_new[9][40];
        llr_in_tmp[9][41]  = llr_new[9][41];
    end
 
    4:begin 
        llr_in_tmp[9][0]  = llr_new[9][0];
        llr_in_tmp[9][1]  = llr_new[9][1];
        llr_in_tmp[9][2]  = llr_new[9][2];
        llr_in_tmp[9][3]  = llr_new[9][3];
        llr_in_tmp[9][4]  = llr_new[9][4];
        llr_in_tmp[9][5]  = llr_new[9][5];
        llr_in_tmp[9][6]  = llr_new[9][6];
        llr_in_tmp[9][7]  = llr_new[9][7];
        llr_in_tmp[9][8]  = llr_new[9][8];
        llr_in_tmp[9][9]  = llr_new[9][9];
        llr_in_tmp[9][10]  = llr_new[9][10];
        llr_in_tmp[9][11]  = llr_new[9][11];
        llr_in_tmp[9][12]  = llr_new[9][12];
        llr_in_tmp[9][13]  = llr_new[9][13];
        llr_in_tmp[9][14]  = llr_new[9][14];
        llr_in_tmp[9][15]  = llr_new[9][15];
        llr_in_tmp[9][16]  = llr_new[9][16];
        llr_in_tmp[9][17]  = llr_new[9][17];
        llr_in_tmp[9][18]  = llr_new[9][18];
        llr_in_tmp[9][19]  = llr_new[9][19];
        llr_in_tmp[9][20]  = llr_new[9][20];
        llr_in_tmp[9][21]  = llr_new[9][21];
        llr_in_tmp[9][22]  = llr_new[9][22];
        llr_in_tmp[9][23]  = llr_new[9][23];
        llr_in_tmp[9][24]  = llr_new[9][24];
        llr_in_tmp[9][25]  = llr_new[9][25];
        llr_in_tmp[9][26]  = llr_new[9][26];
        llr_in_tmp[9][27]  = llr_new[9][27];
        llr_in_tmp[9][28]  = llr_new[9][28];
        llr_in_tmp[9][29]  = llr_new[9][29];
        llr_in_tmp[9][30]  = llr_new[9][30];
        llr_in_tmp[9][31]  = llr_new[9][31];
        llr_in_tmp[9][32]  = llr_new[9][32];
        llr_in_tmp[9][33]  = llr_new[9][33];
        llr_in_tmp[9][34]  = llr_new[9][34];
        llr_in_tmp[9][35]  = llr_new[9][35];
        llr_in_tmp[9][36]  = llr_new[9][36];
        llr_in_tmp[9][37]  = llr_new[9][37];
        llr_in_tmp[9][38]  = llr_new[9][38];
        llr_in_tmp[9][39]  = llr_new[9][39];
        llr_in_tmp[9][40]  = llr_new[9][40];
        llr_in_tmp[9][41]  = llr_new[9][41];
    end
 
    5:begin 
        llr_in_tmp[9][0]  = llr_new[9][28];
        llr_in_tmp[9][1]  = llr_new[9][29];
        llr_in_tmp[9][2]  = llr_new[9][30];
        llr_in_tmp[9][3]  = llr_new[9][31];
        llr_in_tmp[9][4]  = llr_new[9][32];
        llr_in_tmp[9][5]  = llr_new[9][33];
        llr_in_tmp[9][6]  = llr_new[9][34];
        llr_in_tmp[9][7]  = llr_new[9][35];
        llr_in_tmp[9][8]  = llr_new[9][36];
        llr_in_tmp[9][9]  = llr_new[9][37];
        llr_in_tmp[9][10]  = llr_new[9][38];
        llr_in_tmp[9][11]  = llr_new[9][39];
        llr_in_tmp[9][12]  = llr_new[9][40];
        llr_in_tmp[9][13]  = llr_new[9][41];
        llr_in_tmp[9][14]  = llr_new[9][0];
        llr_in_tmp[9][15]  = llr_new[9][1];
        llr_in_tmp[9][16]  = llr_new[9][2];
        llr_in_tmp[9][17]  = llr_new[9][3];
        llr_in_tmp[9][18]  = llr_new[9][4];
        llr_in_tmp[9][19]  = llr_new[9][5];
        llr_in_tmp[9][20]  = llr_new[9][6];
        llr_in_tmp[9][21]  = llr_new[9][7];
        llr_in_tmp[9][22]  = llr_new[9][8];
        llr_in_tmp[9][23]  = llr_new[9][9];
        llr_in_tmp[9][24]  = llr_new[9][10];
        llr_in_tmp[9][25]  = llr_new[9][11];
        llr_in_tmp[9][26]  = llr_new[9][12];
        llr_in_tmp[9][27]  = llr_new[9][13];
        llr_in_tmp[9][28]  = llr_new[9][14];
        llr_in_tmp[9][29]  = llr_new[9][15];
        llr_in_tmp[9][30]  = llr_new[9][16];
        llr_in_tmp[9][31]  = llr_new[9][17];
        llr_in_tmp[9][32]  = llr_new[9][18];
        llr_in_tmp[9][33]  = llr_new[9][19];
        llr_in_tmp[9][34]  = llr_new[9][20];
        llr_in_tmp[9][35]  = llr_new[9][21];
        llr_in_tmp[9][36]  = llr_new[9][22];
        llr_in_tmp[9][37]  = llr_new[9][23];
        llr_in_tmp[9][38]  = llr_new[9][24];
        llr_in_tmp[9][39]  = llr_new[9][25];
        llr_in_tmp[9][40]  = llr_new[9][26];
        llr_in_tmp[9][41]  = llr_new[9][27];
    end
 
    6:begin 
        llr_in_tmp[9][0]  = llr_new[9][0];
        llr_in_tmp[9][1]  = llr_new[9][1];
        llr_in_tmp[9][2]  = llr_new[9][2];
        llr_in_tmp[9][3]  = llr_new[9][3];
        llr_in_tmp[9][4]  = llr_new[9][4];
        llr_in_tmp[9][5]  = llr_new[9][5];
        llr_in_tmp[9][6]  = llr_new[9][6];
        llr_in_tmp[9][7]  = llr_new[9][7];
        llr_in_tmp[9][8]  = llr_new[9][8];
        llr_in_tmp[9][9]  = llr_new[9][9];
        llr_in_tmp[9][10]  = llr_new[9][10];
        llr_in_tmp[9][11]  = llr_new[9][11];
        llr_in_tmp[9][12]  = llr_new[9][12];
        llr_in_tmp[9][13]  = llr_new[9][13];
        llr_in_tmp[9][14]  = llr_new[9][14];
        llr_in_tmp[9][15]  = llr_new[9][15];
        llr_in_tmp[9][16]  = llr_new[9][16];
        llr_in_tmp[9][17]  = llr_new[9][17];
        llr_in_tmp[9][18]  = llr_new[9][18];
        llr_in_tmp[9][19]  = llr_new[9][19];
        llr_in_tmp[9][20]  = llr_new[9][20];
        llr_in_tmp[9][21]  = llr_new[9][21];
        llr_in_tmp[9][22]  = llr_new[9][22];
        llr_in_tmp[9][23]  = llr_new[9][23];
        llr_in_tmp[9][24]  = llr_new[9][24];
        llr_in_tmp[9][25]  = llr_new[9][25];
        llr_in_tmp[9][26]  = llr_new[9][26];
        llr_in_tmp[9][27]  = llr_new[9][27];
        llr_in_tmp[9][28]  = llr_new[9][28];
        llr_in_tmp[9][29]  = llr_new[9][29];
        llr_in_tmp[9][30]  = llr_new[9][30];
        llr_in_tmp[9][31]  = llr_new[9][31];
        llr_in_tmp[9][32]  = llr_new[9][32];
        llr_in_tmp[9][33]  = llr_new[9][33];
        llr_in_tmp[9][34]  = llr_new[9][34];
        llr_in_tmp[9][35]  = llr_new[9][35];
        llr_in_tmp[9][36]  = llr_new[9][36];
        llr_in_tmp[9][37]  = llr_new[9][37];
        llr_in_tmp[9][38]  = llr_new[9][38];
        llr_in_tmp[9][39]  = llr_new[9][39];
        llr_in_tmp[9][40]  = llr_new[9][40];
        llr_in_tmp[9][41]  = llr_new[9][41];
    end
 
    7:begin 
        llr_in_tmp[9][0]  = llr_new[9][0];
        llr_in_tmp[9][1]  = llr_new[9][1];
        llr_in_tmp[9][2]  = llr_new[9][2];
        llr_in_tmp[9][3]  = llr_new[9][3];
        llr_in_tmp[9][4]  = llr_new[9][4];
        llr_in_tmp[9][5]  = llr_new[9][5];
        llr_in_tmp[9][6]  = llr_new[9][6];
        llr_in_tmp[9][7]  = llr_new[9][7];
        llr_in_tmp[9][8]  = llr_new[9][8];
        llr_in_tmp[9][9]  = llr_new[9][9];
        llr_in_tmp[9][10]  = llr_new[9][10];
        llr_in_tmp[9][11]  = llr_new[9][11];
        llr_in_tmp[9][12]  = llr_new[9][12];
        llr_in_tmp[9][13]  = llr_new[9][13];
        llr_in_tmp[9][14]  = llr_new[9][14];
        llr_in_tmp[9][15]  = llr_new[9][15];
        llr_in_tmp[9][16]  = llr_new[9][16];
        llr_in_tmp[9][17]  = llr_new[9][17];
        llr_in_tmp[9][18]  = llr_new[9][18];
        llr_in_tmp[9][19]  = llr_new[9][19];
        llr_in_tmp[9][20]  = llr_new[9][20];
        llr_in_tmp[9][21]  = llr_new[9][21];
        llr_in_tmp[9][22]  = llr_new[9][22];
        llr_in_tmp[9][23]  = llr_new[9][23];
        llr_in_tmp[9][24]  = llr_new[9][24];
        llr_in_tmp[9][25]  = llr_new[9][25];
        llr_in_tmp[9][26]  = llr_new[9][26];
        llr_in_tmp[9][27]  = llr_new[9][27];
        llr_in_tmp[9][28]  = llr_new[9][28];
        llr_in_tmp[9][29]  = llr_new[9][29];
        llr_in_tmp[9][30]  = llr_new[9][30];
        llr_in_tmp[9][31]  = llr_new[9][31];
        llr_in_tmp[9][32]  = llr_new[9][32];
        llr_in_tmp[9][33]  = llr_new[9][33];
        llr_in_tmp[9][34]  = llr_new[9][34];
        llr_in_tmp[9][35]  = llr_new[9][35];
        llr_in_tmp[9][36]  = llr_new[9][36];
        llr_in_tmp[9][37]  = llr_new[9][37];
        llr_in_tmp[9][38]  = llr_new[9][38];
        llr_in_tmp[9][39]  = llr_new[9][39];
        llr_in_tmp[9][40]  = llr_new[9][40];
        llr_in_tmp[9][41]  = llr_new[9][41];
    end
 
endcase
end

if (chk_n_input_valid) begin
case (curr_layer)
    0:begin 
        llr_in_tmp[10][0]  = llr_new[10][0];
        llr_in_tmp[10][1]  = llr_new[10][1];
        llr_in_tmp[10][2]  = llr_new[10][2];
        llr_in_tmp[10][3]  = llr_new[10][3];
        llr_in_tmp[10][4]  = llr_new[10][4];
        llr_in_tmp[10][5]  = llr_new[10][5];
        llr_in_tmp[10][6]  = llr_new[10][6];
        llr_in_tmp[10][7]  = llr_new[10][7];
        llr_in_tmp[10][8]  = llr_new[10][8];
        llr_in_tmp[10][9]  = llr_new[10][9];
        llr_in_tmp[10][10]  = llr_new[10][10];
        llr_in_tmp[10][11]  = llr_new[10][11];
        llr_in_tmp[10][12]  = llr_new[10][12];
        llr_in_tmp[10][13]  = llr_new[10][13];
        llr_in_tmp[10][14]  = llr_new[10][14];
        llr_in_tmp[10][15]  = llr_new[10][15];
        llr_in_tmp[10][16]  = llr_new[10][16];
        llr_in_tmp[10][17]  = llr_new[10][17];
        llr_in_tmp[10][18]  = llr_new[10][18];
        llr_in_tmp[10][19]  = llr_new[10][19];
        llr_in_tmp[10][20]  = llr_new[10][20];
        llr_in_tmp[10][21]  = llr_new[10][21];
        llr_in_tmp[10][22]  = llr_new[10][22];
        llr_in_tmp[10][23]  = llr_new[10][23];
        llr_in_tmp[10][24]  = llr_new[10][24];
        llr_in_tmp[10][25]  = llr_new[10][25];
        llr_in_tmp[10][26]  = llr_new[10][26];
        llr_in_tmp[10][27]  = llr_new[10][27];
        llr_in_tmp[10][28]  = llr_new[10][28];
        llr_in_tmp[10][29]  = llr_new[10][29];
        llr_in_tmp[10][30]  = llr_new[10][30];
        llr_in_tmp[10][31]  = llr_new[10][31];
        llr_in_tmp[10][32]  = llr_new[10][32];
        llr_in_tmp[10][33]  = llr_new[10][33];
        llr_in_tmp[10][34]  = llr_new[10][34];
        llr_in_tmp[10][35]  = llr_new[10][35];
        llr_in_tmp[10][36]  = llr_new[10][36];
        llr_in_tmp[10][37]  = llr_new[10][37];
        llr_in_tmp[10][38]  = llr_new[10][38];
        llr_in_tmp[10][39]  = llr_new[10][39];
        llr_in_tmp[10][40]  = llr_new[10][40];
        llr_in_tmp[10][41]  = llr_new[10][41];
    end
 
    1:begin 
        llr_in_tmp[10][0]  = llr_new[10][0];
        llr_in_tmp[10][1]  = llr_new[10][1];
        llr_in_tmp[10][2]  = llr_new[10][2];
        llr_in_tmp[10][3]  = llr_new[10][3];
        llr_in_tmp[10][4]  = llr_new[10][4];
        llr_in_tmp[10][5]  = llr_new[10][5];
        llr_in_tmp[10][6]  = llr_new[10][6];
        llr_in_tmp[10][7]  = llr_new[10][7];
        llr_in_tmp[10][8]  = llr_new[10][8];
        llr_in_tmp[10][9]  = llr_new[10][9];
        llr_in_tmp[10][10]  = llr_new[10][10];
        llr_in_tmp[10][11]  = llr_new[10][11];
        llr_in_tmp[10][12]  = llr_new[10][12];
        llr_in_tmp[10][13]  = llr_new[10][13];
        llr_in_tmp[10][14]  = llr_new[10][14];
        llr_in_tmp[10][15]  = llr_new[10][15];
        llr_in_tmp[10][16]  = llr_new[10][16];
        llr_in_tmp[10][17]  = llr_new[10][17];
        llr_in_tmp[10][18]  = llr_new[10][18];
        llr_in_tmp[10][19]  = llr_new[10][19];
        llr_in_tmp[10][20]  = llr_new[10][20];
        llr_in_tmp[10][21]  = llr_new[10][21];
        llr_in_tmp[10][22]  = llr_new[10][22];
        llr_in_tmp[10][23]  = llr_new[10][23];
        llr_in_tmp[10][24]  = llr_new[10][24];
        llr_in_tmp[10][25]  = llr_new[10][25];
        llr_in_tmp[10][26]  = llr_new[10][26];
        llr_in_tmp[10][27]  = llr_new[10][27];
        llr_in_tmp[10][28]  = llr_new[10][28];
        llr_in_tmp[10][29]  = llr_new[10][29];
        llr_in_tmp[10][30]  = llr_new[10][30];
        llr_in_tmp[10][31]  = llr_new[10][31];
        llr_in_tmp[10][32]  = llr_new[10][32];
        llr_in_tmp[10][33]  = llr_new[10][33];
        llr_in_tmp[10][34]  = llr_new[10][34];
        llr_in_tmp[10][35]  = llr_new[10][35];
        llr_in_tmp[10][36]  = llr_new[10][36];
        llr_in_tmp[10][37]  = llr_new[10][37];
        llr_in_tmp[10][38]  = llr_new[10][38];
        llr_in_tmp[10][39]  = llr_new[10][39];
        llr_in_tmp[10][40]  = llr_new[10][40];
        llr_in_tmp[10][41]  = llr_new[10][41];
    end
 
    2:begin 
        llr_in_tmp[10][0]  = llr_new[10][41];
        llr_in_tmp[10][1]  = llr_new[10][0];
        llr_in_tmp[10][2]  = llr_new[10][1];
        llr_in_tmp[10][3]  = llr_new[10][2];
        llr_in_tmp[10][4]  = llr_new[10][3];
        llr_in_tmp[10][5]  = llr_new[10][4];
        llr_in_tmp[10][6]  = llr_new[10][5];
        llr_in_tmp[10][7]  = llr_new[10][6];
        llr_in_tmp[10][8]  = llr_new[10][7];
        llr_in_tmp[10][9]  = llr_new[10][8];
        llr_in_tmp[10][10]  = llr_new[10][9];
        llr_in_tmp[10][11]  = llr_new[10][10];
        llr_in_tmp[10][12]  = llr_new[10][11];
        llr_in_tmp[10][13]  = llr_new[10][12];
        llr_in_tmp[10][14]  = llr_new[10][13];
        llr_in_tmp[10][15]  = llr_new[10][14];
        llr_in_tmp[10][16]  = llr_new[10][15];
        llr_in_tmp[10][17]  = llr_new[10][16];
        llr_in_tmp[10][18]  = llr_new[10][17];
        llr_in_tmp[10][19]  = llr_new[10][18];
        llr_in_tmp[10][20]  = llr_new[10][19];
        llr_in_tmp[10][21]  = llr_new[10][20];
        llr_in_tmp[10][22]  = llr_new[10][21];
        llr_in_tmp[10][23]  = llr_new[10][22];
        llr_in_tmp[10][24]  = llr_new[10][23];
        llr_in_tmp[10][25]  = llr_new[10][24];
        llr_in_tmp[10][26]  = llr_new[10][25];
        llr_in_tmp[10][27]  = llr_new[10][26];
        llr_in_tmp[10][28]  = llr_new[10][27];
        llr_in_tmp[10][29]  = llr_new[10][28];
        llr_in_tmp[10][30]  = llr_new[10][29];
        llr_in_tmp[10][31]  = llr_new[10][30];
        llr_in_tmp[10][32]  = llr_new[10][31];
        llr_in_tmp[10][33]  = llr_new[10][32];
        llr_in_tmp[10][34]  = llr_new[10][33];
        llr_in_tmp[10][35]  = llr_new[10][34];
        llr_in_tmp[10][36]  = llr_new[10][35];
        llr_in_tmp[10][37]  = llr_new[10][36];
        llr_in_tmp[10][38]  = llr_new[10][37];
        llr_in_tmp[10][39]  = llr_new[10][38];
        llr_in_tmp[10][40]  = llr_new[10][39];
        llr_in_tmp[10][41]  = llr_new[10][40];
    end
 
    3:begin 
        llr_in_tmp[10][0]  = llr_new[10][15];
        llr_in_tmp[10][1]  = llr_new[10][16];
        llr_in_tmp[10][2]  = llr_new[10][17];
        llr_in_tmp[10][3]  = llr_new[10][18];
        llr_in_tmp[10][4]  = llr_new[10][19];
        llr_in_tmp[10][5]  = llr_new[10][20];
        llr_in_tmp[10][6]  = llr_new[10][21];
        llr_in_tmp[10][7]  = llr_new[10][22];
        llr_in_tmp[10][8]  = llr_new[10][23];
        llr_in_tmp[10][9]  = llr_new[10][24];
        llr_in_tmp[10][10]  = llr_new[10][25];
        llr_in_tmp[10][11]  = llr_new[10][26];
        llr_in_tmp[10][12]  = llr_new[10][27];
        llr_in_tmp[10][13]  = llr_new[10][28];
        llr_in_tmp[10][14]  = llr_new[10][29];
        llr_in_tmp[10][15]  = llr_new[10][30];
        llr_in_tmp[10][16]  = llr_new[10][31];
        llr_in_tmp[10][17]  = llr_new[10][32];
        llr_in_tmp[10][18]  = llr_new[10][33];
        llr_in_tmp[10][19]  = llr_new[10][34];
        llr_in_tmp[10][20]  = llr_new[10][35];
        llr_in_tmp[10][21]  = llr_new[10][36];
        llr_in_tmp[10][22]  = llr_new[10][37];
        llr_in_tmp[10][23]  = llr_new[10][38];
        llr_in_tmp[10][24]  = llr_new[10][39];
        llr_in_tmp[10][25]  = llr_new[10][40];
        llr_in_tmp[10][26]  = llr_new[10][41];
        llr_in_tmp[10][27]  = llr_new[10][0];
        llr_in_tmp[10][28]  = llr_new[10][1];
        llr_in_tmp[10][29]  = llr_new[10][2];
        llr_in_tmp[10][30]  = llr_new[10][3];
        llr_in_tmp[10][31]  = llr_new[10][4];
        llr_in_tmp[10][32]  = llr_new[10][5];
        llr_in_tmp[10][33]  = llr_new[10][6];
        llr_in_tmp[10][34]  = llr_new[10][7];
        llr_in_tmp[10][35]  = llr_new[10][8];
        llr_in_tmp[10][36]  = llr_new[10][9];
        llr_in_tmp[10][37]  = llr_new[10][10];
        llr_in_tmp[10][38]  = llr_new[10][11];
        llr_in_tmp[10][39]  = llr_new[10][12];
        llr_in_tmp[10][40]  = llr_new[10][13];
        llr_in_tmp[10][41]  = llr_new[10][14];
    end
 
    4:begin 
        llr_in_tmp[10][0]  = llr_new[10][0];
        llr_in_tmp[10][1]  = llr_new[10][1];
        llr_in_tmp[10][2]  = llr_new[10][2];
        llr_in_tmp[10][3]  = llr_new[10][3];
        llr_in_tmp[10][4]  = llr_new[10][4];
        llr_in_tmp[10][5]  = llr_new[10][5];
        llr_in_tmp[10][6]  = llr_new[10][6];
        llr_in_tmp[10][7]  = llr_new[10][7];
        llr_in_tmp[10][8]  = llr_new[10][8];
        llr_in_tmp[10][9]  = llr_new[10][9];
        llr_in_tmp[10][10]  = llr_new[10][10];
        llr_in_tmp[10][11]  = llr_new[10][11];
        llr_in_tmp[10][12]  = llr_new[10][12];
        llr_in_tmp[10][13]  = llr_new[10][13];
        llr_in_tmp[10][14]  = llr_new[10][14];
        llr_in_tmp[10][15]  = llr_new[10][15];
        llr_in_tmp[10][16]  = llr_new[10][16];
        llr_in_tmp[10][17]  = llr_new[10][17];
        llr_in_tmp[10][18]  = llr_new[10][18];
        llr_in_tmp[10][19]  = llr_new[10][19];
        llr_in_tmp[10][20]  = llr_new[10][20];
        llr_in_tmp[10][21]  = llr_new[10][21];
        llr_in_tmp[10][22]  = llr_new[10][22];
        llr_in_tmp[10][23]  = llr_new[10][23];
        llr_in_tmp[10][24]  = llr_new[10][24];
        llr_in_tmp[10][25]  = llr_new[10][25];
        llr_in_tmp[10][26]  = llr_new[10][26];
        llr_in_tmp[10][27]  = llr_new[10][27];
        llr_in_tmp[10][28]  = llr_new[10][28];
        llr_in_tmp[10][29]  = llr_new[10][29];
        llr_in_tmp[10][30]  = llr_new[10][30];
        llr_in_tmp[10][31]  = llr_new[10][31];
        llr_in_tmp[10][32]  = llr_new[10][32];
        llr_in_tmp[10][33]  = llr_new[10][33];
        llr_in_tmp[10][34]  = llr_new[10][34];
        llr_in_tmp[10][35]  = llr_new[10][35];
        llr_in_tmp[10][36]  = llr_new[10][36];
        llr_in_tmp[10][37]  = llr_new[10][37];
        llr_in_tmp[10][38]  = llr_new[10][38];
        llr_in_tmp[10][39]  = llr_new[10][39];
        llr_in_tmp[10][40]  = llr_new[10][40];
        llr_in_tmp[10][41]  = llr_new[10][41];
    end
 
    5:begin 
        llr_in_tmp[10][0]  = llr_new[10][0];
        llr_in_tmp[10][1]  = llr_new[10][1];
        llr_in_tmp[10][2]  = llr_new[10][2];
        llr_in_tmp[10][3]  = llr_new[10][3];
        llr_in_tmp[10][4]  = llr_new[10][4];
        llr_in_tmp[10][5]  = llr_new[10][5];
        llr_in_tmp[10][6]  = llr_new[10][6];
        llr_in_tmp[10][7]  = llr_new[10][7];
        llr_in_tmp[10][8]  = llr_new[10][8];
        llr_in_tmp[10][9]  = llr_new[10][9];
        llr_in_tmp[10][10]  = llr_new[10][10];
        llr_in_tmp[10][11]  = llr_new[10][11];
        llr_in_tmp[10][12]  = llr_new[10][12];
        llr_in_tmp[10][13]  = llr_new[10][13];
        llr_in_tmp[10][14]  = llr_new[10][14];
        llr_in_tmp[10][15]  = llr_new[10][15];
        llr_in_tmp[10][16]  = llr_new[10][16];
        llr_in_tmp[10][17]  = llr_new[10][17];
        llr_in_tmp[10][18]  = llr_new[10][18];
        llr_in_tmp[10][19]  = llr_new[10][19];
        llr_in_tmp[10][20]  = llr_new[10][20];
        llr_in_tmp[10][21]  = llr_new[10][21];
        llr_in_tmp[10][22]  = llr_new[10][22];
        llr_in_tmp[10][23]  = llr_new[10][23];
        llr_in_tmp[10][24]  = llr_new[10][24];
        llr_in_tmp[10][25]  = llr_new[10][25];
        llr_in_tmp[10][26]  = llr_new[10][26];
        llr_in_tmp[10][27]  = llr_new[10][27];
        llr_in_tmp[10][28]  = llr_new[10][28];
        llr_in_tmp[10][29]  = llr_new[10][29];
        llr_in_tmp[10][30]  = llr_new[10][30];
        llr_in_tmp[10][31]  = llr_new[10][31];
        llr_in_tmp[10][32]  = llr_new[10][32];
        llr_in_tmp[10][33]  = llr_new[10][33];
        llr_in_tmp[10][34]  = llr_new[10][34];
        llr_in_tmp[10][35]  = llr_new[10][35];
        llr_in_tmp[10][36]  = llr_new[10][36];
        llr_in_tmp[10][37]  = llr_new[10][37];
        llr_in_tmp[10][38]  = llr_new[10][38];
        llr_in_tmp[10][39]  = llr_new[10][39];
        llr_in_tmp[10][40]  = llr_new[10][40];
        llr_in_tmp[10][41]  = llr_new[10][41];
    end
 
    6:begin 
        llr_in_tmp[10][0]  = llr_new[10][12];
        llr_in_tmp[10][1]  = llr_new[10][13];
        llr_in_tmp[10][2]  = llr_new[10][14];
        llr_in_tmp[10][3]  = llr_new[10][15];
        llr_in_tmp[10][4]  = llr_new[10][16];
        llr_in_tmp[10][5]  = llr_new[10][17];
        llr_in_tmp[10][6]  = llr_new[10][18];
        llr_in_tmp[10][7]  = llr_new[10][19];
        llr_in_tmp[10][8]  = llr_new[10][20];
        llr_in_tmp[10][9]  = llr_new[10][21];
        llr_in_tmp[10][10]  = llr_new[10][22];
        llr_in_tmp[10][11]  = llr_new[10][23];
        llr_in_tmp[10][12]  = llr_new[10][24];
        llr_in_tmp[10][13]  = llr_new[10][25];
        llr_in_tmp[10][14]  = llr_new[10][26];
        llr_in_tmp[10][15]  = llr_new[10][27];
        llr_in_tmp[10][16]  = llr_new[10][28];
        llr_in_tmp[10][17]  = llr_new[10][29];
        llr_in_tmp[10][18]  = llr_new[10][30];
        llr_in_tmp[10][19]  = llr_new[10][31];
        llr_in_tmp[10][20]  = llr_new[10][32];
        llr_in_tmp[10][21]  = llr_new[10][33];
        llr_in_tmp[10][22]  = llr_new[10][34];
        llr_in_tmp[10][23]  = llr_new[10][35];
        llr_in_tmp[10][24]  = llr_new[10][36];
        llr_in_tmp[10][25]  = llr_new[10][37];
        llr_in_tmp[10][26]  = llr_new[10][38];
        llr_in_tmp[10][27]  = llr_new[10][39];
        llr_in_tmp[10][28]  = llr_new[10][40];
        llr_in_tmp[10][29]  = llr_new[10][41];
        llr_in_tmp[10][30]  = llr_new[10][0];
        llr_in_tmp[10][31]  = llr_new[10][1];
        llr_in_tmp[10][32]  = llr_new[10][2];
        llr_in_tmp[10][33]  = llr_new[10][3];
        llr_in_tmp[10][34]  = llr_new[10][4];
        llr_in_tmp[10][35]  = llr_new[10][5];
        llr_in_tmp[10][36]  = llr_new[10][6];
        llr_in_tmp[10][37]  = llr_new[10][7];
        llr_in_tmp[10][38]  = llr_new[10][8];
        llr_in_tmp[10][39]  = llr_new[10][9];
        llr_in_tmp[10][40]  = llr_new[10][10];
        llr_in_tmp[10][41]  = llr_new[10][11];
    end
 
    7:begin 
        llr_in_tmp[10][0]  = llr_new[10][0];
        llr_in_tmp[10][1]  = llr_new[10][1];
        llr_in_tmp[10][2]  = llr_new[10][2];
        llr_in_tmp[10][3]  = llr_new[10][3];
        llr_in_tmp[10][4]  = llr_new[10][4];
        llr_in_tmp[10][5]  = llr_new[10][5];
        llr_in_tmp[10][6]  = llr_new[10][6];
        llr_in_tmp[10][7]  = llr_new[10][7];
        llr_in_tmp[10][8]  = llr_new[10][8];
        llr_in_tmp[10][9]  = llr_new[10][9];
        llr_in_tmp[10][10]  = llr_new[10][10];
        llr_in_tmp[10][11]  = llr_new[10][11];
        llr_in_tmp[10][12]  = llr_new[10][12];
        llr_in_tmp[10][13]  = llr_new[10][13];
        llr_in_tmp[10][14]  = llr_new[10][14];
        llr_in_tmp[10][15]  = llr_new[10][15];
        llr_in_tmp[10][16]  = llr_new[10][16];
        llr_in_tmp[10][17]  = llr_new[10][17];
        llr_in_tmp[10][18]  = llr_new[10][18];
        llr_in_tmp[10][19]  = llr_new[10][19];
        llr_in_tmp[10][20]  = llr_new[10][20];
        llr_in_tmp[10][21]  = llr_new[10][21];
        llr_in_tmp[10][22]  = llr_new[10][22];
        llr_in_tmp[10][23]  = llr_new[10][23];
        llr_in_tmp[10][24]  = llr_new[10][24];
        llr_in_tmp[10][25]  = llr_new[10][25];
        llr_in_tmp[10][26]  = llr_new[10][26];
        llr_in_tmp[10][27]  = llr_new[10][27];
        llr_in_tmp[10][28]  = llr_new[10][28];
        llr_in_tmp[10][29]  = llr_new[10][29];
        llr_in_tmp[10][30]  = llr_new[10][30];
        llr_in_tmp[10][31]  = llr_new[10][31];
        llr_in_tmp[10][32]  = llr_new[10][32];
        llr_in_tmp[10][33]  = llr_new[10][33];
        llr_in_tmp[10][34]  = llr_new[10][34];
        llr_in_tmp[10][35]  = llr_new[10][35];
        llr_in_tmp[10][36]  = llr_new[10][36];
        llr_in_tmp[10][37]  = llr_new[10][37];
        llr_in_tmp[10][38]  = llr_new[10][38];
        llr_in_tmp[10][39]  = llr_new[10][39];
        llr_in_tmp[10][40]  = llr_new[10][40];
        llr_in_tmp[10][41]  = llr_new[10][41];
    end
 
endcase
end

if (chk_n_input_valid) begin
case (curr_layer)
    0:begin 
        llr_in_tmp[11][0]  = llr_new[11][0];
        llr_in_tmp[11][1]  = llr_new[11][1];
        llr_in_tmp[11][2]  = llr_new[11][2];
        llr_in_tmp[11][3]  = llr_new[11][3];
        llr_in_tmp[11][4]  = llr_new[11][4];
        llr_in_tmp[11][5]  = llr_new[11][5];
        llr_in_tmp[11][6]  = llr_new[11][6];
        llr_in_tmp[11][7]  = llr_new[11][7];
        llr_in_tmp[11][8]  = llr_new[11][8];
        llr_in_tmp[11][9]  = llr_new[11][9];
        llr_in_tmp[11][10]  = llr_new[11][10];
        llr_in_tmp[11][11]  = llr_new[11][11];
        llr_in_tmp[11][12]  = llr_new[11][12];
        llr_in_tmp[11][13]  = llr_new[11][13];
        llr_in_tmp[11][14]  = llr_new[11][14];
        llr_in_tmp[11][15]  = llr_new[11][15];
        llr_in_tmp[11][16]  = llr_new[11][16];
        llr_in_tmp[11][17]  = llr_new[11][17];
        llr_in_tmp[11][18]  = llr_new[11][18];
        llr_in_tmp[11][19]  = llr_new[11][19];
        llr_in_tmp[11][20]  = llr_new[11][20];
        llr_in_tmp[11][21]  = llr_new[11][21];
        llr_in_tmp[11][22]  = llr_new[11][22];
        llr_in_tmp[11][23]  = llr_new[11][23];
        llr_in_tmp[11][24]  = llr_new[11][24];
        llr_in_tmp[11][25]  = llr_new[11][25];
        llr_in_tmp[11][26]  = llr_new[11][26];
        llr_in_tmp[11][27]  = llr_new[11][27];
        llr_in_tmp[11][28]  = llr_new[11][28];
        llr_in_tmp[11][29]  = llr_new[11][29];
        llr_in_tmp[11][30]  = llr_new[11][30];
        llr_in_tmp[11][31]  = llr_new[11][31];
        llr_in_tmp[11][32]  = llr_new[11][32];
        llr_in_tmp[11][33]  = llr_new[11][33];
        llr_in_tmp[11][34]  = llr_new[11][34];
        llr_in_tmp[11][35]  = llr_new[11][35];
        llr_in_tmp[11][36]  = llr_new[11][36];
        llr_in_tmp[11][37]  = llr_new[11][37];
        llr_in_tmp[11][38]  = llr_new[11][38];
        llr_in_tmp[11][39]  = llr_new[11][39];
        llr_in_tmp[11][40]  = llr_new[11][40];
        llr_in_tmp[11][41]  = llr_new[11][41];
    end
 
    1:begin 
        llr_in_tmp[11][0]  = llr_new[11][0];
        llr_in_tmp[11][1]  = llr_new[11][1];
        llr_in_tmp[11][2]  = llr_new[11][2];
        llr_in_tmp[11][3]  = llr_new[11][3];
        llr_in_tmp[11][4]  = llr_new[11][4];
        llr_in_tmp[11][5]  = llr_new[11][5];
        llr_in_tmp[11][6]  = llr_new[11][6];
        llr_in_tmp[11][7]  = llr_new[11][7];
        llr_in_tmp[11][8]  = llr_new[11][8];
        llr_in_tmp[11][9]  = llr_new[11][9];
        llr_in_tmp[11][10]  = llr_new[11][10];
        llr_in_tmp[11][11]  = llr_new[11][11];
        llr_in_tmp[11][12]  = llr_new[11][12];
        llr_in_tmp[11][13]  = llr_new[11][13];
        llr_in_tmp[11][14]  = llr_new[11][14];
        llr_in_tmp[11][15]  = llr_new[11][15];
        llr_in_tmp[11][16]  = llr_new[11][16];
        llr_in_tmp[11][17]  = llr_new[11][17];
        llr_in_tmp[11][18]  = llr_new[11][18];
        llr_in_tmp[11][19]  = llr_new[11][19];
        llr_in_tmp[11][20]  = llr_new[11][20];
        llr_in_tmp[11][21]  = llr_new[11][21];
        llr_in_tmp[11][22]  = llr_new[11][22];
        llr_in_tmp[11][23]  = llr_new[11][23];
        llr_in_tmp[11][24]  = llr_new[11][24];
        llr_in_tmp[11][25]  = llr_new[11][25];
        llr_in_tmp[11][26]  = llr_new[11][26];
        llr_in_tmp[11][27]  = llr_new[11][27];
        llr_in_tmp[11][28]  = llr_new[11][28];
        llr_in_tmp[11][29]  = llr_new[11][29];
        llr_in_tmp[11][30]  = llr_new[11][30];
        llr_in_tmp[11][31]  = llr_new[11][31];
        llr_in_tmp[11][32]  = llr_new[11][32];
        llr_in_tmp[11][33]  = llr_new[11][33];
        llr_in_tmp[11][34]  = llr_new[11][34];
        llr_in_tmp[11][35]  = llr_new[11][35];
        llr_in_tmp[11][36]  = llr_new[11][36];
        llr_in_tmp[11][37]  = llr_new[11][37];
        llr_in_tmp[11][38]  = llr_new[11][38];
        llr_in_tmp[11][39]  = llr_new[11][39];
        llr_in_tmp[11][40]  = llr_new[11][40];
        llr_in_tmp[11][41]  = llr_new[11][41];
    end
 
    2:begin 
        llr_in_tmp[11][0]  = llr_new[11][0];
        llr_in_tmp[11][1]  = llr_new[11][1];
        llr_in_tmp[11][2]  = llr_new[11][2];
        llr_in_tmp[11][3]  = llr_new[11][3];
        llr_in_tmp[11][4]  = llr_new[11][4];
        llr_in_tmp[11][5]  = llr_new[11][5];
        llr_in_tmp[11][6]  = llr_new[11][6];
        llr_in_tmp[11][7]  = llr_new[11][7];
        llr_in_tmp[11][8]  = llr_new[11][8];
        llr_in_tmp[11][9]  = llr_new[11][9];
        llr_in_tmp[11][10]  = llr_new[11][10];
        llr_in_tmp[11][11]  = llr_new[11][11];
        llr_in_tmp[11][12]  = llr_new[11][12];
        llr_in_tmp[11][13]  = llr_new[11][13];
        llr_in_tmp[11][14]  = llr_new[11][14];
        llr_in_tmp[11][15]  = llr_new[11][15];
        llr_in_tmp[11][16]  = llr_new[11][16];
        llr_in_tmp[11][17]  = llr_new[11][17];
        llr_in_tmp[11][18]  = llr_new[11][18];
        llr_in_tmp[11][19]  = llr_new[11][19];
        llr_in_tmp[11][20]  = llr_new[11][20];
        llr_in_tmp[11][21]  = llr_new[11][21];
        llr_in_tmp[11][22]  = llr_new[11][22];
        llr_in_tmp[11][23]  = llr_new[11][23];
        llr_in_tmp[11][24]  = llr_new[11][24];
        llr_in_tmp[11][25]  = llr_new[11][25];
        llr_in_tmp[11][26]  = llr_new[11][26];
        llr_in_tmp[11][27]  = llr_new[11][27];
        llr_in_tmp[11][28]  = llr_new[11][28];
        llr_in_tmp[11][29]  = llr_new[11][29];
        llr_in_tmp[11][30]  = llr_new[11][30];
        llr_in_tmp[11][31]  = llr_new[11][31];
        llr_in_tmp[11][32]  = llr_new[11][32];
        llr_in_tmp[11][33]  = llr_new[11][33];
        llr_in_tmp[11][34]  = llr_new[11][34];
        llr_in_tmp[11][35]  = llr_new[11][35];
        llr_in_tmp[11][36]  = llr_new[11][36];
        llr_in_tmp[11][37]  = llr_new[11][37];
        llr_in_tmp[11][38]  = llr_new[11][38];
        llr_in_tmp[11][39]  = llr_new[11][39];
        llr_in_tmp[11][40]  = llr_new[11][40];
        llr_in_tmp[11][41]  = llr_new[11][41];
    end
 
    3:begin 
        llr_in_tmp[11][0]  = llr_new[11][6];
        llr_in_tmp[11][1]  = llr_new[11][7];
        llr_in_tmp[11][2]  = llr_new[11][8];
        llr_in_tmp[11][3]  = llr_new[11][9];
        llr_in_tmp[11][4]  = llr_new[11][10];
        llr_in_tmp[11][5]  = llr_new[11][11];
        llr_in_tmp[11][6]  = llr_new[11][12];
        llr_in_tmp[11][7]  = llr_new[11][13];
        llr_in_tmp[11][8]  = llr_new[11][14];
        llr_in_tmp[11][9]  = llr_new[11][15];
        llr_in_tmp[11][10]  = llr_new[11][16];
        llr_in_tmp[11][11]  = llr_new[11][17];
        llr_in_tmp[11][12]  = llr_new[11][18];
        llr_in_tmp[11][13]  = llr_new[11][19];
        llr_in_tmp[11][14]  = llr_new[11][20];
        llr_in_tmp[11][15]  = llr_new[11][21];
        llr_in_tmp[11][16]  = llr_new[11][22];
        llr_in_tmp[11][17]  = llr_new[11][23];
        llr_in_tmp[11][18]  = llr_new[11][24];
        llr_in_tmp[11][19]  = llr_new[11][25];
        llr_in_tmp[11][20]  = llr_new[11][26];
        llr_in_tmp[11][21]  = llr_new[11][27];
        llr_in_tmp[11][22]  = llr_new[11][28];
        llr_in_tmp[11][23]  = llr_new[11][29];
        llr_in_tmp[11][24]  = llr_new[11][30];
        llr_in_tmp[11][25]  = llr_new[11][31];
        llr_in_tmp[11][26]  = llr_new[11][32];
        llr_in_tmp[11][27]  = llr_new[11][33];
        llr_in_tmp[11][28]  = llr_new[11][34];
        llr_in_tmp[11][29]  = llr_new[11][35];
        llr_in_tmp[11][30]  = llr_new[11][36];
        llr_in_tmp[11][31]  = llr_new[11][37];
        llr_in_tmp[11][32]  = llr_new[11][38];
        llr_in_tmp[11][33]  = llr_new[11][39];
        llr_in_tmp[11][34]  = llr_new[11][40];
        llr_in_tmp[11][35]  = llr_new[11][41];
        llr_in_tmp[11][36]  = llr_new[11][0];
        llr_in_tmp[11][37]  = llr_new[11][1];
        llr_in_tmp[11][38]  = llr_new[11][2];
        llr_in_tmp[11][39]  = llr_new[11][3];
        llr_in_tmp[11][40]  = llr_new[11][4];
        llr_in_tmp[11][41]  = llr_new[11][5];
    end
 
    4:begin 
        llr_in_tmp[11][0]  = llr_new[11][3];
        llr_in_tmp[11][1]  = llr_new[11][4];
        llr_in_tmp[11][2]  = llr_new[11][5];
        llr_in_tmp[11][3]  = llr_new[11][6];
        llr_in_tmp[11][4]  = llr_new[11][7];
        llr_in_tmp[11][5]  = llr_new[11][8];
        llr_in_tmp[11][6]  = llr_new[11][9];
        llr_in_tmp[11][7]  = llr_new[11][10];
        llr_in_tmp[11][8]  = llr_new[11][11];
        llr_in_tmp[11][9]  = llr_new[11][12];
        llr_in_tmp[11][10]  = llr_new[11][13];
        llr_in_tmp[11][11]  = llr_new[11][14];
        llr_in_tmp[11][12]  = llr_new[11][15];
        llr_in_tmp[11][13]  = llr_new[11][16];
        llr_in_tmp[11][14]  = llr_new[11][17];
        llr_in_tmp[11][15]  = llr_new[11][18];
        llr_in_tmp[11][16]  = llr_new[11][19];
        llr_in_tmp[11][17]  = llr_new[11][20];
        llr_in_tmp[11][18]  = llr_new[11][21];
        llr_in_tmp[11][19]  = llr_new[11][22];
        llr_in_tmp[11][20]  = llr_new[11][23];
        llr_in_tmp[11][21]  = llr_new[11][24];
        llr_in_tmp[11][22]  = llr_new[11][25];
        llr_in_tmp[11][23]  = llr_new[11][26];
        llr_in_tmp[11][24]  = llr_new[11][27];
        llr_in_tmp[11][25]  = llr_new[11][28];
        llr_in_tmp[11][26]  = llr_new[11][29];
        llr_in_tmp[11][27]  = llr_new[11][30];
        llr_in_tmp[11][28]  = llr_new[11][31];
        llr_in_tmp[11][29]  = llr_new[11][32];
        llr_in_tmp[11][30]  = llr_new[11][33];
        llr_in_tmp[11][31]  = llr_new[11][34];
        llr_in_tmp[11][32]  = llr_new[11][35];
        llr_in_tmp[11][33]  = llr_new[11][36];
        llr_in_tmp[11][34]  = llr_new[11][37];
        llr_in_tmp[11][35]  = llr_new[11][38];
        llr_in_tmp[11][36]  = llr_new[11][39];
        llr_in_tmp[11][37]  = llr_new[11][40];
        llr_in_tmp[11][38]  = llr_new[11][41];
        llr_in_tmp[11][39]  = llr_new[11][0];
        llr_in_tmp[11][40]  = llr_new[11][1];
        llr_in_tmp[11][41]  = llr_new[11][2];
    end
 
    5:begin 
        llr_in_tmp[11][0]  = llr_new[11][27];
        llr_in_tmp[11][1]  = llr_new[11][28];
        llr_in_tmp[11][2]  = llr_new[11][29];
        llr_in_tmp[11][3]  = llr_new[11][30];
        llr_in_tmp[11][4]  = llr_new[11][31];
        llr_in_tmp[11][5]  = llr_new[11][32];
        llr_in_tmp[11][6]  = llr_new[11][33];
        llr_in_tmp[11][7]  = llr_new[11][34];
        llr_in_tmp[11][8]  = llr_new[11][35];
        llr_in_tmp[11][9]  = llr_new[11][36];
        llr_in_tmp[11][10]  = llr_new[11][37];
        llr_in_tmp[11][11]  = llr_new[11][38];
        llr_in_tmp[11][12]  = llr_new[11][39];
        llr_in_tmp[11][13]  = llr_new[11][40];
        llr_in_tmp[11][14]  = llr_new[11][41];
        llr_in_tmp[11][15]  = llr_new[11][0];
        llr_in_tmp[11][16]  = llr_new[11][1];
        llr_in_tmp[11][17]  = llr_new[11][2];
        llr_in_tmp[11][18]  = llr_new[11][3];
        llr_in_tmp[11][19]  = llr_new[11][4];
        llr_in_tmp[11][20]  = llr_new[11][5];
        llr_in_tmp[11][21]  = llr_new[11][6];
        llr_in_tmp[11][22]  = llr_new[11][7];
        llr_in_tmp[11][23]  = llr_new[11][8];
        llr_in_tmp[11][24]  = llr_new[11][9];
        llr_in_tmp[11][25]  = llr_new[11][10];
        llr_in_tmp[11][26]  = llr_new[11][11];
        llr_in_tmp[11][27]  = llr_new[11][12];
        llr_in_tmp[11][28]  = llr_new[11][13];
        llr_in_tmp[11][29]  = llr_new[11][14];
        llr_in_tmp[11][30]  = llr_new[11][15];
        llr_in_tmp[11][31]  = llr_new[11][16];
        llr_in_tmp[11][32]  = llr_new[11][17];
        llr_in_tmp[11][33]  = llr_new[11][18];
        llr_in_tmp[11][34]  = llr_new[11][19];
        llr_in_tmp[11][35]  = llr_new[11][20];
        llr_in_tmp[11][36]  = llr_new[11][21];
        llr_in_tmp[11][37]  = llr_new[11][22];
        llr_in_tmp[11][38]  = llr_new[11][23];
        llr_in_tmp[11][39]  = llr_new[11][24];
        llr_in_tmp[11][40]  = llr_new[11][25];
        llr_in_tmp[11][41]  = llr_new[11][26];
    end
 
    6:begin 
        llr_in_tmp[11][0]  = llr_new[11][0];
        llr_in_tmp[11][1]  = llr_new[11][1];
        llr_in_tmp[11][2]  = llr_new[11][2];
        llr_in_tmp[11][3]  = llr_new[11][3];
        llr_in_tmp[11][4]  = llr_new[11][4];
        llr_in_tmp[11][5]  = llr_new[11][5];
        llr_in_tmp[11][6]  = llr_new[11][6];
        llr_in_tmp[11][7]  = llr_new[11][7];
        llr_in_tmp[11][8]  = llr_new[11][8];
        llr_in_tmp[11][9]  = llr_new[11][9];
        llr_in_tmp[11][10]  = llr_new[11][10];
        llr_in_tmp[11][11]  = llr_new[11][11];
        llr_in_tmp[11][12]  = llr_new[11][12];
        llr_in_tmp[11][13]  = llr_new[11][13];
        llr_in_tmp[11][14]  = llr_new[11][14];
        llr_in_tmp[11][15]  = llr_new[11][15];
        llr_in_tmp[11][16]  = llr_new[11][16];
        llr_in_tmp[11][17]  = llr_new[11][17];
        llr_in_tmp[11][18]  = llr_new[11][18];
        llr_in_tmp[11][19]  = llr_new[11][19];
        llr_in_tmp[11][20]  = llr_new[11][20];
        llr_in_tmp[11][21]  = llr_new[11][21];
        llr_in_tmp[11][22]  = llr_new[11][22];
        llr_in_tmp[11][23]  = llr_new[11][23];
        llr_in_tmp[11][24]  = llr_new[11][24];
        llr_in_tmp[11][25]  = llr_new[11][25];
        llr_in_tmp[11][26]  = llr_new[11][26];
        llr_in_tmp[11][27]  = llr_new[11][27];
        llr_in_tmp[11][28]  = llr_new[11][28];
        llr_in_tmp[11][29]  = llr_new[11][29];
        llr_in_tmp[11][30]  = llr_new[11][30];
        llr_in_tmp[11][31]  = llr_new[11][31];
        llr_in_tmp[11][32]  = llr_new[11][32];
        llr_in_tmp[11][33]  = llr_new[11][33];
        llr_in_tmp[11][34]  = llr_new[11][34];
        llr_in_tmp[11][35]  = llr_new[11][35];
        llr_in_tmp[11][36]  = llr_new[11][36];
        llr_in_tmp[11][37]  = llr_new[11][37];
        llr_in_tmp[11][38]  = llr_new[11][38];
        llr_in_tmp[11][39]  = llr_new[11][39];
        llr_in_tmp[11][40]  = llr_new[11][40];
        llr_in_tmp[11][41]  = llr_new[11][41];
    end
 
    7:begin 
        llr_in_tmp[11][0]  = llr_new[11][0];
        llr_in_tmp[11][1]  = llr_new[11][1];
        llr_in_tmp[11][2]  = llr_new[11][2];
        llr_in_tmp[11][3]  = llr_new[11][3];
        llr_in_tmp[11][4]  = llr_new[11][4];
        llr_in_tmp[11][5]  = llr_new[11][5];
        llr_in_tmp[11][6]  = llr_new[11][6];
        llr_in_tmp[11][7]  = llr_new[11][7];
        llr_in_tmp[11][8]  = llr_new[11][8];
        llr_in_tmp[11][9]  = llr_new[11][9];
        llr_in_tmp[11][10]  = llr_new[11][10];
        llr_in_tmp[11][11]  = llr_new[11][11];
        llr_in_tmp[11][12]  = llr_new[11][12];
        llr_in_tmp[11][13]  = llr_new[11][13];
        llr_in_tmp[11][14]  = llr_new[11][14];
        llr_in_tmp[11][15]  = llr_new[11][15];
        llr_in_tmp[11][16]  = llr_new[11][16];
        llr_in_tmp[11][17]  = llr_new[11][17];
        llr_in_tmp[11][18]  = llr_new[11][18];
        llr_in_tmp[11][19]  = llr_new[11][19];
        llr_in_tmp[11][20]  = llr_new[11][20];
        llr_in_tmp[11][21]  = llr_new[11][21];
        llr_in_tmp[11][22]  = llr_new[11][22];
        llr_in_tmp[11][23]  = llr_new[11][23];
        llr_in_tmp[11][24]  = llr_new[11][24];
        llr_in_tmp[11][25]  = llr_new[11][25];
        llr_in_tmp[11][26]  = llr_new[11][26];
        llr_in_tmp[11][27]  = llr_new[11][27];
        llr_in_tmp[11][28]  = llr_new[11][28];
        llr_in_tmp[11][29]  = llr_new[11][29];
        llr_in_tmp[11][30]  = llr_new[11][30];
        llr_in_tmp[11][31]  = llr_new[11][31];
        llr_in_tmp[11][32]  = llr_new[11][32];
        llr_in_tmp[11][33]  = llr_new[11][33];
        llr_in_tmp[11][34]  = llr_new[11][34];
        llr_in_tmp[11][35]  = llr_new[11][35];
        llr_in_tmp[11][36]  = llr_new[11][36];
        llr_in_tmp[11][37]  = llr_new[11][37];
        llr_in_tmp[11][38]  = llr_new[11][38];
        llr_in_tmp[11][39]  = llr_new[11][39];
        llr_in_tmp[11][40]  = llr_new[11][40];
        llr_in_tmp[11][41]  = llr_new[11][41];
    end
 
endcase
end

if (chk_n_input_valid) begin
case (curr_layer)
    0:begin 
        llr_in_tmp[12][0]  = llr_new[12][0];
        llr_in_tmp[12][1]  = llr_new[12][1];
        llr_in_tmp[12][2]  = llr_new[12][2];
        llr_in_tmp[12][3]  = llr_new[12][3];
        llr_in_tmp[12][4]  = llr_new[12][4];
        llr_in_tmp[12][5]  = llr_new[12][5];
        llr_in_tmp[12][6]  = llr_new[12][6];
        llr_in_tmp[12][7]  = llr_new[12][7];
        llr_in_tmp[12][8]  = llr_new[12][8];
        llr_in_tmp[12][9]  = llr_new[12][9];
        llr_in_tmp[12][10]  = llr_new[12][10];
        llr_in_tmp[12][11]  = llr_new[12][11];
        llr_in_tmp[12][12]  = llr_new[12][12];
        llr_in_tmp[12][13]  = llr_new[12][13];
        llr_in_tmp[12][14]  = llr_new[12][14];
        llr_in_tmp[12][15]  = llr_new[12][15];
        llr_in_tmp[12][16]  = llr_new[12][16];
        llr_in_tmp[12][17]  = llr_new[12][17];
        llr_in_tmp[12][18]  = llr_new[12][18];
        llr_in_tmp[12][19]  = llr_new[12][19];
        llr_in_tmp[12][20]  = llr_new[12][20];
        llr_in_tmp[12][21]  = llr_new[12][21];
        llr_in_tmp[12][22]  = llr_new[12][22];
        llr_in_tmp[12][23]  = llr_new[12][23];
        llr_in_tmp[12][24]  = llr_new[12][24];
        llr_in_tmp[12][25]  = llr_new[12][25];
        llr_in_tmp[12][26]  = llr_new[12][26];
        llr_in_tmp[12][27]  = llr_new[12][27];
        llr_in_tmp[12][28]  = llr_new[12][28];
        llr_in_tmp[12][29]  = llr_new[12][29];
        llr_in_tmp[12][30]  = llr_new[12][30];
        llr_in_tmp[12][31]  = llr_new[12][31];
        llr_in_tmp[12][32]  = llr_new[12][32];
        llr_in_tmp[12][33]  = llr_new[12][33];
        llr_in_tmp[12][34]  = llr_new[12][34];
        llr_in_tmp[12][35]  = llr_new[12][35];
        llr_in_tmp[12][36]  = llr_new[12][36];
        llr_in_tmp[12][37]  = llr_new[12][37];
        llr_in_tmp[12][38]  = llr_new[12][38];
        llr_in_tmp[12][39]  = llr_new[12][39];
        llr_in_tmp[12][40]  = llr_new[12][40];
        llr_in_tmp[12][41]  = llr_new[12][41];
    end
 
    1:begin 
        llr_in_tmp[12][0]  = llr_new[12][0];
        llr_in_tmp[12][1]  = llr_new[12][1];
        llr_in_tmp[12][2]  = llr_new[12][2];
        llr_in_tmp[12][3]  = llr_new[12][3];
        llr_in_tmp[12][4]  = llr_new[12][4];
        llr_in_tmp[12][5]  = llr_new[12][5];
        llr_in_tmp[12][6]  = llr_new[12][6];
        llr_in_tmp[12][7]  = llr_new[12][7];
        llr_in_tmp[12][8]  = llr_new[12][8];
        llr_in_tmp[12][9]  = llr_new[12][9];
        llr_in_tmp[12][10]  = llr_new[12][10];
        llr_in_tmp[12][11]  = llr_new[12][11];
        llr_in_tmp[12][12]  = llr_new[12][12];
        llr_in_tmp[12][13]  = llr_new[12][13];
        llr_in_tmp[12][14]  = llr_new[12][14];
        llr_in_tmp[12][15]  = llr_new[12][15];
        llr_in_tmp[12][16]  = llr_new[12][16];
        llr_in_tmp[12][17]  = llr_new[12][17];
        llr_in_tmp[12][18]  = llr_new[12][18];
        llr_in_tmp[12][19]  = llr_new[12][19];
        llr_in_tmp[12][20]  = llr_new[12][20];
        llr_in_tmp[12][21]  = llr_new[12][21];
        llr_in_tmp[12][22]  = llr_new[12][22];
        llr_in_tmp[12][23]  = llr_new[12][23];
        llr_in_tmp[12][24]  = llr_new[12][24];
        llr_in_tmp[12][25]  = llr_new[12][25];
        llr_in_tmp[12][26]  = llr_new[12][26];
        llr_in_tmp[12][27]  = llr_new[12][27];
        llr_in_tmp[12][28]  = llr_new[12][28];
        llr_in_tmp[12][29]  = llr_new[12][29];
        llr_in_tmp[12][30]  = llr_new[12][30];
        llr_in_tmp[12][31]  = llr_new[12][31];
        llr_in_tmp[12][32]  = llr_new[12][32];
        llr_in_tmp[12][33]  = llr_new[12][33];
        llr_in_tmp[12][34]  = llr_new[12][34];
        llr_in_tmp[12][35]  = llr_new[12][35];
        llr_in_tmp[12][36]  = llr_new[12][36];
        llr_in_tmp[12][37]  = llr_new[12][37];
        llr_in_tmp[12][38]  = llr_new[12][38];
        llr_in_tmp[12][39]  = llr_new[12][39];
        llr_in_tmp[12][40]  = llr_new[12][40];
        llr_in_tmp[12][41]  = llr_new[12][41];
    end
 
    2:begin 
        llr_in_tmp[12][0]  = llr_new[12][0];
        llr_in_tmp[12][1]  = llr_new[12][1];
        llr_in_tmp[12][2]  = llr_new[12][2];
        llr_in_tmp[12][3]  = llr_new[12][3];
        llr_in_tmp[12][4]  = llr_new[12][4];
        llr_in_tmp[12][5]  = llr_new[12][5];
        llr_in_tmp[12][6]  = llr_new[12][6];
        llr_in_tmp[12][7]  = llr_new[12][7];
        llr_in_tmp[12][8]  = llr_new[12][8];
        llr_in_tmp[12][9]  = llr_new[12][9];
        llr_in_tmp[12][10]  = llr_new[12][10];
        llr_in_tmp[12][11]  = llr_new[12][11];
        llr_in_tmp[12][12]  = llr_new[12][12];
        llr_in_tmp[12][13]  = llr_new[12][13];
        llr_in_tmp[12][14]  = llr_new[12][14];
        llr_in_tmp[12][15]  = llr_new[12][15];
        llr_in_tmp[12][16]  = llr_new[12][16];
        llr_in_tmp[12][17]  = llr_new[12][17];
        llr_in_tmp[12][18]  = llr_new[12][18];
        llr_in_tmp[12][19]  = llr_new[12][19];
        llr_in_tmp[12][20]  = llr_new[12][20];
        llr_in_tmp[12][21]  = llr_new[12][21];
        llr_in_tmp[12][22]  = llr_new[12][22];
        llr_in_tmp[12][23]  = llr_new[12][23];
        llr_in_tmp[12][24]  = llr_new[12][24];
        llr_in_tmp[12][25]  = llr_new[12][25];
        llr_in_tmp[12][26]  = llr_new[12][26];
        llr_in_tmp[12][27]  = llr_new[12][27];
        llr_in_tmp[12][28]  = llr_new[12][28];
        llr_in_tmp[12][29]  = llr_new[12][29];
        llr_in_tmp[12][30]  = llr_new[12][30];
        llr_in_tmp[12][31]  = llr_new[12][31];
        llr_in_tmp[12][32]  = llr_new[12][32];
        llr_in_tmp[12][33]  = llr_new[12][33];
        llr_in_tmp[12][34]  = llr_new[12][34];
        llr_in_tmp[12][35]  = llr_new[12][35];
        llr_in_tmp[12][36]  = llr_new[12][36];
        llr_in_tmp[12][37]  = llr_new[12][37];
        llr_in_tmp[12][38]  = llr_new[12][38];
        llr_in_tmp[12][39]  = llr_new[12][39];
        llr_in_tmp[12][40]  = llr_new[12][40];
        llr_in_tmp[12][41]  = llr_new[12][41];
    end
 
    3:begin 
        llr_in_tmp[12][0]  = llr_new[12][0];
        llr_in_tmp[12][1]  = llr_new[12][1];
        llr_in_tmp[12][2]  = llr_new[12][2];
        llr_in_tmp[12][3]  = llr_new[12][3];
        llr_in_tmp[12][4]  = llr_new[12][4];
        llr_in_tmp[12][5]  = llr_new[12][5];
        llr_in_tmp[12][6]  = llr_new[12][6];
        llr_in_tmp[12][7]  = llr_new[12][7];
        llr_in_tmp[12][8]  = llr_new[12][8];
        llr_in_tmp[12][9]  = llr_new[12][9];
        llr_in_tmp[12][10]  = llr_new[12][10];
        llr_in_tmp[12][11]  = llr_new[12][11];
        llr_in_tmp[12][12]  = llr_new[12][12];
        llr_in_tmp[12][13]  = llr_new[12][13];
        llr_in_tmp[12][14]  = llr_new[12][14];
        llr_in_tmp[12][15]  = llr_new[12][15];
        llr_in_tmp[12][16]  = llr_new[12][16];
        llr_in_tmp[12][17]  = llr_new[12][17];
        llr_in_tmp[12][18]  = llr_new[12][18];
        llr_in_tmp[12][19]  = llr_new[12][19];
        llr_in_tmp[12][20]  = llr_new[12][20];
        llr_in_tmp[12][21]  = llr_new[12][21];
        llr_in_tmp[12][22]  = llr_new[12][22];
        llr_in_tmp[12][23]  = llr_new[12][23];
        llr_in_tmp[12][24]  = llr_new[12][24];
        llr_in_tmp[12][25]  = llr_new[12][25];
        llr_in_tmp[12][26]  = llr_new[12][26];
        llr_in_tmp[12][27]  = llr_new[12][27];
        llr_in_tmp[12][28]  = llr_new[12][28];
        llr_in_tmp[12][29]  = llr_new[12][29];
        llr_in_tmp[12][30]  = llr_new[12][30];
        llr_in_tmp[12][31]  = llr_new[12][31];
        llr_in_tmp[12][32]  = llr_new[12][32];
        llr_in_tmp[12][33]  = llr_new[12][33];
        llr_in_tmp[12][34]  = llr_new[12][34];
        llr_in_tmp[12][35]  = llr_new[12][35];
        llr_in_tmp[12][36]  = llr_new[12][36];
        llr_in_tmp[12][37]  = llr_new[12][37];
        llr_in_tmp[12][38]  = llr_new[12][38];
        llr_in_tmp[12][39]  = llr_new[12][39];
        llr_in_tmp[12][40]  = llr_new[12][40];
        llr_in_tmp[12][41]  = llr_new[12][41];
    end
 
    4:begin 
        llr_in_tmp[12][0]  = llr_new[12][28];
        llr_in_tmp[12][1]  = llr_new[12][29];
        llr_in_tmp[12][2]  = llr_new[12][30];
        llr_in_tmp[12][3]  = llr_new[12][31];
        llr_in_tmp[12][4]  = llr_new[12][32];
        llr_in_tmp[12][5]  = llr_new[12][33];
        llr_in_tmp[12][6]  = llr_new[12][34];
        llr_in_tmp[12][7]  = llr_new[12][35];
        llr_in_tmp[12][8]  = llr_new[12][36];
        llr_in_tmp[12][9]  = llr_new[12][37];
        llr_in_tmp[12][10]  = llr_new[12][38];
        llr_in_tmp[12][11]  = llr_new[12][39];
        llr_in_tmp[12][12]  = llr_new[12][40];
        llr_in_tmp[12][13]  = llr_new[12][41];
        llr_in_tmp[12][14]  = llr_new[12][0];
        llr_in_tmp[12][15]  = llr_new[12][1];
        llr_in_tmp[12][16]  = llr_new[12][2];
        llr_in_tmp[12][17]  = llr_new[12][3];
        llr_in_tmp[12][18]  = llr_new[12][4];
        llr_in_tmp[12][19]  = llr_new[12][5];
        llr_in_tmp[12][20]  = llr_new[12][6];
        llr_in_tmp[12][21]  = llr_new[12][7];
        llr_in_tmp[12][22]  = llr_new[12][8];
        llr_in_tmp[12][23]  = llr_new[12][9];
        llr_in_tmp[12][24]  = llr_new[12][10];
        llr_in_tmp[12][25]  = llr_new[12][11];
        llr_in_tmp[12][26]  = llr_new[12][12];
        llr_in_tmp[12][27]  = llr_new[12][13];
        llr_in_tmp[12][28]  = llr_new[12][14];
        llr_in_tmp[12][29]  = llr_new[12][15];
        llr_in_tmp[12][30]  = llr_new[12][16];
        llr_in_tmp[12][31]  = llr_new[12][17];
        llr_in_tmp[12][32]  = llr_new[12][18];
        llr_in_tmp[12][33]  = llr_new[12][19];
        llr_in_tmp[12][34]  = llr_new[12][20];
        llr_in_tmp[12][35]  = llr_new[12][21];
        llr_in_tmp[12][36]  = llr_new[12][22];
        llr_in_tmp[12][37]  = llr_new[12][23];
        llr_in_tmp[12][38]  = llr_new[12][24];
        llr_in_tmp[12][39]  = llr_new[12][25];
        llr_in_tmp[12][40]  = llr_new[12][26];
        llr_in_tmp[12][41]  = llr_new[12][27];
    end
 
    5:begin 
        llr_in_tmp[12][0]  = llr_new[12][0];
        llr_in_tmp[12][1]  = llr_new[12][1];
        llr_in_tmp[12][2]  = llr_new[12][2];
        llr_in_tmp[12][3]  = llr_new[12][3];
        llr_in_tmp[12][4]  = llr_new[12][4];
        llr_in_tmp[12][5]  = llr_new[12][5];
        llr_in_tmp[12][6]  = llr_new[12][6];
        llr_in_tmp[12][7]  = llr_new[12][7];
        llr_in_tmp[12][8]  = llr_new[12][8];
        llr_in_tmp[12][9]  = llr_new[12][9];
        llr_in_tmp[12][10]  = llr_new[12][10];
        llr_in_tmp[12][11]  = llr_new[12][11];
        llr_in_tmp[12][12]  = llr_new[12][12];
        llr_in_tmp[12][13]  = llr_new[12][13];
        llr_in_tmp[12][14]  = llr_new[12][14];
        llr_in_tmp[12][15]  = llr_new[12][15];
        llr_in_tmp[12][16]  = llr_new[12][16];
        llr_in_tmp[12][17]  = llr_new[12][17];
        llr_in_tmp[12][18]  = llr_new[12][18];
        llr_in_tmp[12][19]  = llr_new[12][19];
        llr_in_tmp[12][20]  = llr_new[12][20];
        llr_in_tmp[12][21]  = llr_new[12][21];
        llr_in_tmp[12][22]  = llr_new[12][22];
        llr_in_tmp[12][23]  = llr_new[12][23];
        llr_in_tmp[12][24]  = llr_new[12][24];
        llr_in_tmp[12][25]  = llr_new[12][25];
        llr_in_tmp[12][26]  = llr_new[12][26];
        llr_in_tmp[12][27]  = llr_new[12][27];
        llr_in_tmp[12][28]  = llr_new[12][28];
        llr_in_tmp[12][29]  = llr_new[12][29];
        llr_in_tmp[12][30]  = llr_new[12][30];
        llr_in_tmp[12][31]  = llr_new[12][31];
        llr_in_tmp[12][32]  = llr_new[12][32];
        llr_in_tmp[12][33]  = llr_new[12][33];
        llr_in_tmp[12][34]  = llr_new[12][34];
        llr_in_tmp[12][35]  = llr_new[12][35];
        llr_in_tmp[12][36]  = llr_new[12][36];
        llr_in_tmp[12][37]  = llr_new[12][37];
        llr_in_tmp[12][38]  = llr_new[12][38];
        llr_in_tmp[12][39]  = llr_new[12][39];
        llr_in_tmp[12][40]  = llr_new[12][40];
        llr_in_tmp[12][41]  = llr_new[12][41];
    end
 
    6:begin 
        llr_in_tmp[12][0]  = llr_new[12][0];
        llr_in_tmp[12][1]  = llr_new[12][1];
        llr_in_tmp[12][2]  = llr_new[12][2];
        llr_in_tmp[12][3]  = llr_new[12][3];
        llr_in_tmp[12][4]  = llr_new[12][4];
        llr_in_tmp[12][5]  = llr_new[12][5];
        llr_in_tmp[12][6]  = llr_new[12][6];
        llr_in_tmp[12][7]  = llr_new[12][7];
        llr_in_tmp[12][8]  = llr_new[12][8];
        llr_in_tmp[12][9]  = llr_new[12][9];
        llr_in_tmp[12][10]  = llr_new[12][10];
        llr_in_tmp[12][11]  = llr_new[12][11];
        llr_in_tmp[12][12]  = llr_new[12][12];
        llr_in_tmp[12][13]  = llr_new[12][13];
        llr_in_tmp[12][14]  = llr_new[12][14];
        llr_in_tmp[12][15]  = llr_new[12][15];
        llr_in_tmp[12][16]  = llr_new[12][16];
        llr_in_tmp[12][17]  = llr_new[12][17];
        llr_in_tmp[12][18]  = llr_new[12][18];
        llr_in_tmp[12][19]  = llr_new[12][19];
        llr_in_tmp[12][20]  = llr_new[12][20];
        llr_in_tmp[12][21]  = llr_new[12][21];
        llr_in_tmp[12][22]  = llr_new[12][22];
        llr_in_tmp[12][23]  = llr_new[12][23];
        llr_in_tmp[12][24]  = llr_new[12][24];
        llr_in_tmp[12][25]  = llr_new[12][25];
        llr_in_tmp[12][26]  = llr_new[12][26];
        llr_in_tmp[12][27]  = llr_new[12][27];
        llr_in_tmp[12][28]  = llr_new[12][28];
        llr_in_tmp[12][29]  = llr_new[12][29];
        llr_in_tmp[12][30]  = llr_new[12][30];
        llr_in_tmp[12][31]  = llr_new[12][31];
        llr_in_tmp[12][32]  = llr_new[12][32];
        llr_in_tmp[12][33]  = llr_new[12][33];
        llr_in_tmp[12][34]  = llr_new[12][34];
        llr_in_tmp[12][35]  = llr_new[12][35];
        llr_in_tmp[12][36]  = llr_new[12][36];
        llr_in_tmp[12][37]  = llr_new[12][37];
        llr_in_tmp[12][38]  = llr_new[12][38];
        llr_in_tmp[12][39]  = llr_new[12][39];
        llr_in_tmp[12][40]  = llr_new[12][40];
        llr_in_tmp[12][41]  = llr_new[12][41];
    end
 
    7:begin 
        llr_in_tmp[12][0]  = llr_new[12][13];
        llr_in_tmp[12][1]  = llr_new[12][14];
        llr_in_tmp[12][2]  = llr_new[12][15];
        llr_in_tmp[12][3]  = llr_new[12][16];
        llr_in_tmp[12][4]  = llr_new[12][17];
        llr_in_tmp[12][5]  = llr_new[12][18];
        llr_in_tmp[12][6]  = llr_new[12][19];
        llr_in_tmp[12][7]  = llr_new[12][20];
        llr_in_tmp[12][8]  = llr_new[12][21];
        llr_in_tmp[12][9]  = llr_new[12][22];
        llr_in_tmp[12][10]  = llr_new[12][23];
        llr_in_tmp[12][11]  = llr_new[12][24];
        llr_in_tmp[12][12]  = llr_new[12][25];
        llr_in_tmp[12][13]  = llr_new[12][26];
        llr_in_tmp[12][14]  = llr_new[12][27];
        llr_in_tmp[12][15]  = llr_new[12][28];
        llr_in_tmp[12][16]  = llr_new[12][29];
        llr_in_tmp[12][17]  = llr_new[12][30];
        llr_in_tmp[12][18]  = llr_new[12][31];
        llr_in_tmp[12][19]  = llr_new[12][32];
        llr_in_tmp[12][20]  = llr_new[12][33];
        llr_in_tmp[12][21]  = llr_new[12][34];
        llr_in_tmp[12][22]  = llr_new[12][35];
        llr_in_tmp[12][23]  = llr_new[12][36];
        llr_in_tmp[12][24]  = llr_new[12][37];
        llr_in_tmp[12][25]  = llr_new[12][38];
        llr_in_tmp[12][26]  = llr_new[12][39];
        llr_in_tmp[12][27]  = llr_new[12][40];
        llr_in_tmp[12][28]  = llr_new[12][41];
        llr_in_tmp[12][29]  = llr_new[12][0];
        llr_in_tmp[12][30]  = llr_new[12][1];
        llr_in_tmp[12][31]  = llr_new[12][2];
        llr_in_tmp[12][32]  = llr_new[12][3];
        llr_in_tmp[12][33]  = llr_new[12][4];
        llr_in_tmp[12][34]  = llr_new[12][5];
        llr_in_tmp[12][35]  = llr_new[12][6];
        llr_in_tmp[12][36]  = llr_new[12][7];
        llr_in_tmp[12][37]  = llr_new[12][8];
        llr_in_tmp[12][38]  = llr_new[12][9];
        llr_in_tmp[12][39]  = llr_new[12][10];
        llr_in_tmp[12][40]  = llr_new[12][11];
        llr_in_tmp[12][41]  = llr_new[12][12];
    end
 
endcase
end

if (chk_n_input_valid) begin
case (curr_layer)
    0:begin 
        llr_in_tmp[13][0]  = llr_new[13][0];
        llr_in_tmp[13][1]  = llr_new[13][1];
        llr_in_tmp[13][2]  = llr_new[13][2];
        llr_in_tmp[13][3]  = llr_new[13][3];
        llr_in_tmp[13][4]  = llr_new[13][4];
        llr_in_tmp[13][5]  = llr_new[13][5];
        llr_in_tmp[13][6]  = llr_new[13][6];
        llr_in_tmp[13][7]  = llr_new[13][7];
        llr_in_tmp[13][8]  = llr_new[13][8];
        llr_in_tmp[13][9]  = llr_new[13][9];
        llr_in_tmp[13][10]  = llr_new[13][10];
        llr_in_tmp[13][11]  = llr_new[13][11];
        llr_in_tmp[13][12]  = llr_new[13][12];
        llr_in_tmp[13][13]  = llr_new[13][13];
        llr_in_tmp[13][14]  = llr_new[13][14];
        llr_in_tmp[13][15]  = llr_new[13][15];
        llr_in_tmp[13][16]  = llr_new[13][16];
        llr_in_tmp[13][17]  = llr_new[13][17];
        llr_in_tmp[13][18]  = llr_new[13][18];
        llr_in_tmp[13][19]  = llr_new[13][19];
        llr_in_tmp[13][20]  = llr_new[13][20];
        llr_in_tmp[13][21]  = llr_new[13][21];
        llr_in_tmp[13][22]  = llr_new[13][22];
        llr_in_tmp[13][23]  = llr_new[13][23];
        llr_in_tmp[13][24]  = llr_new[13][24];
        llr_in_tmp[13][25]  = llr_new[13][25];
        llr_in_tmp[13][26]  = llr_new[13][26];
        llr_in_tmp[13][27]  = llr_new[13][27];
        llr_in_tmp[13][28]  = llr_new[13][28];
        llr_in_tmp[13][29]  = llr_new[13][29];
        llr_in_tmp[13][30]  = llr_new[13][30];
        llr_in_tmp[13][31]  = llr_new[13][31];
        llr_in_tmp[13][32]  = llr_new[13][32];
        llr_in_tmp[13][33]  = llr_new[13][33];
        llr_in_tmp[13][34]  = llr_new[13][34];
        llr_in_tmp[13][35]  = llr_new[13][35];
        llr_in_tmp[13][36]  = llr_new[13][36];
        llr_in_tmp[13][37]  = llr_new[13][37];
        llr_in_tmp[13][38]  = llr_new[13][38];
        llr_in_tmp[13][39]  = llr_new[13][39];
        llr_in_tmp[13][40]  = llr_new[13][40];
        llr_in_tmp[13][41]  = llr_new[13][41];
    end
 
    1:begin 
        llr_in_tmp[13][0]  = llr_new[13][0];
        llr_in_tmp[13][1]  = llr_new[13][1];
        llr_in_tmp[13][2]  = llr_new[13][2];
        llr_in_tmp[13][3]  = llr_new[13][3];
        llr_in_tmp[13][4]  = llr_new[13][4];
        llr_in_tmp[13][5]  = llr_new[13][5];
        llr_in_tmp[13][6]  = llr_new[13][6];
        llr_in_tmp[13][7]  = llr_new[13][7];
        llr_in_tmp[13][8]  = llr_new[13][8];
        llr_in_tmp[13][9]  = llr_new[13][9];
        llr_in_tmp[13][10]  = llr_new[13][10];
        llr_in_tmp[13][11]  = llr_new[13][11];
        llr_in_tmp[13][12]  = llr_new[13][12];
        llr_in_tmp[13][13]  = llr_new[13][13];
        llr_in_tmp[13][14]  = llr_new[13][14];
        llr_in_tmp[13][15]  = llr_new[13][15];
        llr_in_tmp[13][16]  = llr_new[13][16];
        llr_in_tmp[13][17]  = llr_new[13][17];
        llr_in_tmp[13][18]  = llr_new[13][18];
        llr_in_tmp[13][19]  = llr_new[13][19];
        llr_in_tmp[13][20]  = llr_new[13][20];
        llr_in_tmp[13][21]  = llr_new[13][21];
        llr_in_tmp[13][22]  = llr_new[13][22];
        llr_in_tmp[13][23]  = llr_new[13][23];
        llr_in_tmp[13][24]  = llr_new[13][24];
        llr_in_tmp[13][25]  = llr_new[13][25];
        llr_in_tmp[13][26]  = llr_new[13][26];
        llr_in_tmp[13][27]  = llr_new[13][27];
        llr_in_tmp[13][28]  = llr_new[13][28];
        llr_in_tmp[13][29]  = llr_new[13][29];
        llr_in_tmp[13][30]  = llr_new[13][30];
        llr_in_tmp[13][31]  = llr_new[13][31];
        llr_in_tmp[13][32]  = llr_new[13][32];
        llr_in_tmp[13][33]  = llr_new[13][33];
        llr_in_tmp[13][34]  = llr_new[13][34];
        llr_in_tmp[13][35]  = llr_new[13][35];
        llr_in_tmp[13][36]  = llr_new[13][36];
        llr_in_tmp[13][37]  = llr_new[13][37];
        llr_in_tmp[13][38]  = llr_new[13][38];
        llr_in_tmp[13][39]  = llr_new[13][39];
        llr_in_tmp[13][40]  = llr_new[13][40];
        llr_in_tmp[13][41]  = llr_new[13][41];
    end
 
    2:begin 
        llr_in_tmp[13][0]  = llr_new[13][0];
        llr_in_tmp[13][1]  = llr_new[13][1];
        llr_in_tmp[13][2]  = llr_new[13][2];
        llr_in_tmp[13][3]  = llr_new[13][3];
        llr_in_tmp[13][4]  = llr_new[13][4];
        llr_in_tmp[13][5]  = llr_new[13][5];
        llr_in_tmp[13][6]  = llr_new[13][6];
        llr_in_tmp[13][7]  = llr_new[13][7];
        llr_in_tmp[13][8]  = llr_new[13][8];
        llr_in_tmp[13][9]  = llr_new[13][9];
        llr_in_tmp[13][10]  = llr_new[13][10];
        llr_in_tmp[13][11]  = llr_new[13][11];
        llr_in_tmp[13][12]  = llr_new[13][12];
        llr_in_tmp[13][13]  = llr_new[13][13];
        llr_in_tmp[13][14]  = llr_new[13][14];
        llr_in_tmp[13][15]  = llr_new[13][15];
        llr_in_tmp[13][16]  = llr_new[13][16];
        llr_in_tmp[13][17]  = llr_new[13][17];
        llr_in_tmp[13][18]  = llr_new[13][18];
        llr_in_tmp[13][19]  = llr_new[13][19];
        llr_in_tmp[13][20]  = llr_new[13][20];
        llr_in_tmp[13][21]  = llr_new[13][21];
        llr_in_tmp[13][22]  = llr_new[13][22];
        llr_in_tmp[13][23]  = llr_new[13][23];
        llr_in_tmp[13][24]  = llr_new[13][24];
        llr_in_tmp[13][25]  = llr_new[13][25];
        llr_in_tmp[13][26]  = llr_new[13][26];
        llr_in_tmp[13][27]  = llr_new[13][27];
        llr_in_tmp[13][28]  = llr_new[13][28];
        llr_in_tmp[13][29]  = llr_new[13][29];
        llr_in_tmp[13][30]  = llr_new[13][30];
        llr_in_tmp[13][31]  = llr_new[13][31];
        llr_in_tmp[13][32]  = llr_new[13][32];
        llr_in_tmp[13][33]  = llr_new[13][33];
        llr_in_tmp[13][34]  = llr_new[13][34];
        llr_in_tmp[13][35]  = llr_new[13][35];
        llr_in_tmp[13][36]  = llr_new[13][36];
        llr_in_tmp[13][37]  = llr_new[13][37];
        llr_in_tmp[13][38]  = llr_new[13][38];
        llr_in_tmp[13][39]  = llr_new[13][39];
        llr_in_tmp[13][40]  = llr_new[13][40];
        llr_in_tmp[13][41]  = llr_new[13][41];
    end
 
    3:begin 
        llr_in_tmp[13][0]  = llr_new[13][0];
        llr_in_tmp[13][1]  = llr_new[13][1];
        llr_in_tmp[13][2]  = llr_new[13][2];
        llr_in_tmp[13][3]  = llr_new[13][3];
        llr_in_tmp[13][4]  = llr_new[13][4];
        llr_in_tmp[13][5]  = llr_new[13][5];
        llr_in_tmp[13][6]  = llr_new[13][6];
        llr_in_tmp[13][7]  = llr_new[13][7];
        llr_in_tmp[13][8]  = llr_new[13][8];
        llr_in_tmp[13][9]  = llr_new[13][9];
        llr_in_tmp[13][10]  = llr_new[13][10];
        llr_in_tmp[13][11]  = llr_new[13][11];
        llr_in_tmp[13][12]  = llr_new[13][12];
        llr_in_tmp[13][13]  = llr_new[13][13];
        llr_in_tmp[13][14]  = llr_new[13][14];
        llr_in_tmp[13][15]  = llr_new[13][15];
        llr_in_tmp[13][16]  = llr_new[13][16];
        llr_in_tmp[13][17]  = llr_new[13][17];
        llr_in_tmp[13][18]  = llr_new[13][18];
        llr_in_tmp[13][19]  = llr_new[13][19];
        llr_in_tmp[13][20]  = llr_new[13][20];
        llr_in_tmp[13][21]  = llr_new[13][21];
        llr_in_tmp[13][22]  = llr_new[13][22];
        llr_in_tmp[13][23]  = llr_new[13][23];
        llr_in_tmp[13][24]  = llr_new[13][24];
        llr_in_tmp[13][25]  = llr_new[13][25];
        llr_in_tmp[13][26]  = llr_new[13][26];
        llr_in_tmp[13][27]  = llr_new[13][27];
        llr_in_tmp[13][28]  = llr_new[13][28];
        llr_in_tmp[13][29]  = llr_new[13][29];
        llr_in_tmp[13][30]  = llr_new[13][30];
        llr_in_tmp[13][31]  = llr_new[13][31];
        llr_in_tmp[13][32]  = llr_new[13][32];
        llr_in_tmp[13][33]  = llr_new[13][33];
        llr_in_tmp[13][34]  = llr_new[13][34];
        llr_in_tmp[13][35]  = llr_new[13][35];
        llr_in_tmp[13][36]  = llr_new[13][36];
        llr_in_tmp[13][37]  = llr_new[13][37];
        llr_in_tmp[13][38]  = llr_new[13][38];
        llr_in_tmp[13][39]  = llr_new[13][39];
        llr_in_tmp[13][40]  = llr_new[13][40];
        llr_in_tmp[13][41]  = llr_new[13][41];
    end
 
    4:begin 
        llr_in_tmp[13][0]  = llr_new[13][0];
        llr_in_tmp[13][1]  = llr_new[13][1];
        llr_in_tmp[13][2]  = llr_new[13][2];
        llr_in_tmp[13][3]  = llr_new[13][3];
        llr_in_tmp[13][4]  = llr_new[13][4];
        llr_in_tmp[13][5]  = llr_new[13][5];
        llr_in_tmp[13][6]  = llr_new[13][6];
        llr_in_tmp[13][7]  = llr_new[13][7];
        llr_in_tmp[13][8]  = llr_new[13][8];
        llr_in_tmp[13][9]  = llr_new[13][9];
        llr_in_tmp[13][10]  = llr_new[13][10];
        llr_in_tmp[13][11]  = llr_new[13][11];
        llr_in_tmp[13][12]  = llr_new[13][12];
        llr_in_tmp[13][13]  = llr_new[13][13];
        llr_in_tmp[13][14]  = llr_new[13][14];
        llr_in_tmp[13][15]  = llr_new[13][15];
        llr_in_tmp[13][16]  = llr_new[13][16];
        llr_in_tmp[13][17]  = llr_new[13][17];
        llr_in_tmp[13][18]  = llr_new[13][18];
        llr_in_tmp[13][19]  = llr_new[13][19];
        llr_in_tmp[13][20]  = llr_new[13][20];
        llr_in_tmp[13][21]  = llr_new[13][21];
        llr_in_tmp[13][22]  = llr_new[13][22];
        llr_in_tmp[13][23]  = llr_new[13][23];
        llr_in_tmp[13][24]  = llr_new[13][24];
        llr_in_tmp[13][25]  = llr_new[13][25];
        llr_in_tmp[13][26]  = llr_new[13][26];
        llr_in_tmp[13][27]  = llr_new[13][27];
        llr_in_tmp[13][28]  = llr_new[13][28];
        llr_in_tmp[13][29]  = llr_new[13][29];
        llr_in_tmp[13][30]  = llr_new[13][30];
        llr_in_tmp[13][31]  = llr_new[13][31];
        llr_in_tmp[13][32]  = llr_new[13][32];
        llr_in_tmp[13][33]  = llr_new[13][33];
        llr_in_tmp[13][34]  = llr_new[13][34];
        llr_in_tmp[13][35]  = llr_new[13][35];
        llr_in_tmp[13][36]  = llr_new[13][36];
        llr_in_tmp[13][37]  = llr_new[13][37];
        llr_in_tmp[13][38]  = llr_new[13][38];
        llr_in_tmp[13][39]  = llr_new[13][39];
        llr_in_tmp[13][40]  = llr_new[13][40];
        llr_in_tmp[13][41]  = llr_new[13][41];
    end
 
    5:begin 
        llr_in_tmp[13][0]  = llr_new[13][23];
        llr_in_tmp[13][1]  = llr_new[13][24];
        llr_in_tmp[13][2]  = llr_new[13][25];
        llr_in_tmp[13][3]  = llr_new[13][26];
        llr_in_tmp[13][4]  = llr_new[13][27];
        llr_in_tmp[13][5]  = llr_new[13][28];
        llr_in_tmp[13][6]  = llr_new[13][29];
        llr_in_tmp[13][7]  = llr_new[13][30];
        llr_in_tmp[13][8]  = llr_new[13][31];
        llr_in_tmp[13][9]  = llr_new[13][32];
        llr_in_tmp[13][10]  = llr_new[13][33];
        llr_in_tmp[13][11]  = llr_new[13][34];
        llr_in_tmp[13][12]  = llr_new[13][35];
        llr_in_tmp[13][13]  = llr_new[13][36];
        llr_in_tmp[13][14]  = llr_new[13][37];
        llr_in_tmp[13][15]  = llr_new[13][38];
        llr_in_tmp[13][16]  = llr_new[13][39];
        llr_in_tmp[13][17]  = llr_new[13][40];
        llr_in_tmp[13][18]  = llr_new[13][41];
        llr_in_tmp[13][19]  = llr_new[13][0];
        llr_in_tmp[13][20]  = llr_new[13][1];
        llr_in_tmp[13][21]  = llr_new[13][2];
        llr_in_tmp[13][22]  = llr_new[13][3];
        llr_in_tmp[13][23]  = llr_new[13][4];
        llr_in_tmp[13][24]  = llr_new[13][5];
        llr_in_tmp[13][25]  = llr_new[13][6];
        llr_in_tmp[13][26]  = llr_new[13][7];
        llr_in_tmp[13][27]  = llr_new[13][8];
        llr_in_tmp[13][28]  = llr_new[13][9];
        llr_in_tmp[13][29]  = llr_new[13][10];
        llr_in_tmp[13][30]  = llr_new[13][11];
        llr_in_tmp[13][31]  = llr_new[13][12];
        llr_in_tmp[13][32]  = llr_new[13][13];
        llr_in_tmp[13][33]  = llr_new[13][14];
        llr_in_tmp[13][34]  = llr_new[13][15];
        llr_in_tmp[13][35]  = llr_new[13][16];
        llr_in_tmp[13][36]  = llr_new[13][17];
        llr_in_tmp[13][37]  = llr_new[13][18];
        llr_in_tmp[13][38]  = llr_new[13][19];
        llr_in_tmp[13][39]  = llr_new[13][20];
        llr_in_tmp[13][40]  = llr_new[13][21];
        llr_in_tmp[13][41]  = llr_new[13][22];
    end
 
    6:begin 
        llr_in_tmp[13][0]  = llr_new[13][0];
        llr_in_tmp[13][1]  = llr_new[13][1];
        llr_in_tmp[13][2]  = llr_new[13][2];
        llr_in_tmp[13][3]  = llr_new[13][3];
        llr_in_tmp[13][4]  = llr_new[13][4];
        llr_in_tmp[13][5]  = llr_new[13][5];
        llr_in_tmp[13][6]  = llr_new[13][6];
        llr_in_tmp[13][7]  = llr_new[13][7];
        llr_in_tmp[13][8]  = llr_new[13][8];
        llr_in_tmp[13][9]  = llr_new[13][9];
        llr_in_tmp[13][10]  = llr_new[13][10];
        llr_in_tmp[13][11]  = llr_new[13][11];
        llr_in_tmp[13][12]  = llr_new[13][12];
        llr_in_tmp[13][13]  = llr_new[13][13];
        llr_in_tmp[13][14]  = llr_new[13][14];
        llr_in_tmp[13][15]  = llr_new[13][15];
        llr_in_tmp[13][16]  = llr_new[13][16];
        llr_in_tmp[13][17]  = llr_new[13][17];
        llr_in_tmp[13][18]  = llr_new[13][18];
        llr_in_tmp[13][19]  = llr_new[13][19];
        llr_in_tmp[13][20]  = llr_new[13][20];
        llr_in_tmp[13][21]  = llr_new[13][21];
        llr_in_tmp[13][22]  = llr_new[13][22];
        llr_in_tmp[13][23]  = llr_new[13][23];
        llr_in_tmp[13][24]  = llr_new[13][24];
        llr_in_tmp[13][25]  = llr_new[13][25];
        llr_in_tmp[13][26]  = llr_new[13][26];
        llr_in_tmp[13][27]  = llr_new[13][27];
        llr_in_tmp[13][28]  = llr_new[13][28];
        llr_in_tmp[13][29]  = llr_new[13][29];
        llr_in_tmp[13][30]  = llr_new[13][30];
        llr_in_tmp[13][31]  = llr_new[13][31];
        llr_in_tmp[13][32]  = llr_new[13][32];
        llr_in_tmp[13][33]  = llr_new[13][33];
        llr_in_tmp[13][34]  = llr_new[13][34];
        llr_in_tmp[13][35]  = llr_new[13][35];
        llr_in_tmp[13][36]  = llr_new[13][36];
        llr_in_tmp[13][37]  = llr_new[13][37];
        llr_in_tmp[13][38]  = llr_new[13][38];
        llr_in_tmp[13][39]  = llr_new[13][39];
        llr_in_tmp[13][40]  = llr_new[13][40];
        llr_in_tmp[13][41]  = llr_new[13][41];
    end
 
    7:begin 
        llr_in_tmp[13][0]  = llr_new[13][0];
        llr_in_tmp[13][1]  = llr_new[13][1];
        llr_in_tmp[13][2]  = llr_new[13][2];
        llr_in_tmp[13][3]  = llr_new[13][3];
        llr_in_tmp[13][4]  = llr_new[13][4];
        llr_in_tmp[13][5]  = llr_new[13][5];
        llr_in_tmp[13][6]  = llr_new[13][6];
        llr_in_tmp[13][7]  = llr_new[13][7];
        llr_in_tmp[13][8]  = llr_new[13][8];
        llr_in_tmp[13][9]  = llr_new[13][9];
        llr_in_tmp[13][10]  = llr_new[13][10];
        llr_in_tmp[13][11]  = llr_new[13][11];
        llr_in_tmp[13][12]  = llr_new[13][12];
        llr_in_tmp[13][13]  = llr_new[13][13];
        llr_in_tmp[13][14]  = llr_new[13][14];
        llr_in_tmp[13][15]  = llr_new[13][15];
        llr_in_tmp[13][16]  = llr_new[13][16];
        llr_in_tmp[13][17]  = llr_new[13][17];
        llr_in_tmp[13][18]  = llr_new[13][18];
        llr_in_tmp[13][19]  = llr_new[13][19];
        llr_in_tmp[13][20]  = llr_new[13][20];
        llr_in_tmp[13][21]  = llr_new[13][21];
        llr_in_tmp[13][22]  = llr_new[13][22];
        llr_in_tmp[13][23]  = llr_new[13][23];
        llr_in_tmp[13][24]  = llr_new[13][24];
        llr_in_tmp[13][25]  = llr_new[13][25];
        llr_in_tmp[13][26]  = llr_new[13][26];
        llr_in_tmp[13][27]  = llr_new[13][27];
        llr_in_tmp[13][28]  = llr_new[13][28];
        llr_in_tmp[13][29]  = llr_new[13][29];
        llr_in_tmp[13][30]  = llr_new[13][30];
        llr_in_tmp[13][31]  = llr_new[13][31];
        llr_in_tmp[13][32]  = llr_new[13][32];
        llr_in_tmp[13][33]  = llr_new[13][33];
        llr_in_tmp[13][34]  = llr_new[13][34];
        llr_in_tmp[13][35]  = llr_new[13][35];
        llr_in_tmp[13][36]  = llr_new[13][36];
        llr_in_tmp[13][37]  = llr_new[13][37];
        llr_in_tmp[13][38]  = llr_new[13][38];
        llr_in_tmp[13][39]  = llr_new[13][39];
        llr_in_tmp[13][40]  = llr_new[13][40];
        llr_in_tmp[13][41]  = llr_new[13][41];
    end
 
endcase
end

if (chk_n_input_valid) begin
case (curr_layer)
    0:begin 
        llr_in_tmp[14][0]  = llr_new[14][0];
        llr_in_tmp[14][1]  = llr_new[14][1];
        llr_in_tmp[14][2]  = llr_new[14][2];
        llr_in_tmp[14][3]  = llr_new[14][3];
        llr_in_tmp[14][4]  = llr_new[14][4];
        llr_in_tmp[14][5]  = llr_new[14][5];
        llr_in_tmp[14][6]  = llr_new[14][6];
        llr_in_tmp[14][7]  = llr_new[14][7];
        llr_in_tmp[14][8]  = llr_new[14][8];
        llr_in_tmp[14][9]  = llr_new[14][9];
        llr_in_tmp[14][10]  = llr_new[14][10];
        llr_in_tmp[14][11]  = llr_new[14][11];
        llr_in_tmp[14][12]  = llr_new[14][12];
        llr_in_tmp[14][13]  = llr_new[14][13];
        llr_in_tmp[14][14]  = llr_new[14][14];
        llr_in_tmp[14][15]  = llr_new[14][15];
        llr_in_tmp[14][16]  = llr_new[14][16];
        llr_in_tmp[14][17]  = llr_new[14][17];
        llr_in_tmp[14][18]  = llr_new[14][18];
        llr_in_tmp[14][19]  = llr_new[14][19];
        llr_in_tmp[14][20]  = llr_new[14][20];
        llr_in_tmp[14][21]  = llr_new[14][21];
        llr_in_tmp[14][22]  = llr_new[14][22];
        llr_in_tmp[14][23]  = llr_new[14][23];
        llr_in_tmp[14][24]  = llr_new[14][24];
        llr_in_tmp[14][25]  = llr_new[14][25];
        llr_in_tmp[14][26]  = llr_new[14][26];
        llr_in_tmp[14][27]  = llr_new[14][27];
        llr_in_tmp[14][28]  = llr_new[14][28];
        llr_in_tmp[14][29]  = llr_new[14][29];
        llr_in_tmp[14][30]  = llr_new[14][30];
        llr_in_tmp[14][31]  = llr_new[14][31];
        llr_in_tmp[14][32]  = llr_new[14][32];
        llr_in_tmp[14][33]  = llr_new[14][33];
        llr_in_tmp[14][34]  = llr_new[14][34];
        llr_in_tmp[14][35]  = llr_new[14][35];
        llr_in_tmp[14][36]  = llr_new[14][36];
        llr_in_tmp[14][37]  = llr_new[14][37];
        llr_in_tmp[14][38]  = llr_new[14][38];
        llr_in_tmp[14][39]  = llr_new[14][39];
        llr_in_tmp[14][40]  = llr_new[14][40];
        llr_in_tmp[14][41]  = llr_new[14][41];
    end
 
    1:begin 
        llr_in_tmp[14][0]  = llr_new[14][0];
        llr_in_tmp[14][1]  = llr_new[14][1];
        llr_in_tmp[14][2]  = llr_new[14][2];
        llr_in_tmp[14][3]  = llr_new[14][3];
        llr_in_tmp[14][4]  = llr_new[14][4];
        llr_in_tmp[14][5]  = llr_new[14][5];
        llr_in_tmp[14][6]  = llr_new[14][6];
        llr_in_tmp[14][7]  = llr_new[14][7];
        llr_in_tmp[14][8]  = llr_new[14][8];
        llr_in_tmp[14][9]  = llr_new[14][9];
        llr_in_tmp[14][10]  = llr_new[14][10];
        llr_in_tmp[14][11]  = llr_new[14][11];
        llr_in_tmp[14][12]  = llr_new[14][12];
        llr_in_tmp[14][13]  = llr_new[14][13];
        llr_in_tmp[14][14]  = llr_new[14][14];
        llr_in_tmp[14][15]  = llr_new[14][15];
        llr_in_tmp[14][16]  = llr_new[14][16];
        llr_in_tmp[14][17]  = llr_new[14][17];
        llr_in_tmp[14][18]  = llr_new[14][18];
        llr_in_tmp[14][19]  = llr_new[14][19];
        llr_in_tmp[14][20]  = llr_new[14][20];
        llr_in_tmp[14][21]  = llr_new[14][21];
        llr_in_tmp[14][22]  = llr_new[14][22];
        llr_in_tmp[14][23]  = llr_new[14][23];
        llr_in_tmp[14][24]  = llr_new[14][24];
        llr_in_tmp[14][25]  = llr_new[14][25];
        llr_in_tmp[14][26]  = llr_new[14][26];
        llr_in_tmp[14][27]  = llr_new[14][27];
        llr_in_tmp[14][28]  = llr_new[14][28];
        llr_in_tmp[14][29]  = llr_new[14][29];
        llr_in_tmp[14][30]  = llr_new[14][30];
        llr_in_tmp[14][31]  = llr_new[14][31];
        llr_in_tmp[14][32]  = llr_new[14][32];
        llr_in_tmp[14][33]  = llr_new[14][33];
        llr_in_tmp[14][34]  = llr_new[14][34];
        llr_in_tmp[14][35]  = llr_new[14][35];
        llr_in_tmp[14][36]  = llr_new[14][36];
        llr_in_tmp[14][37]  = llr_new[14][37];
        llr_in_tmp[14][38]  = llr_new[14][38];
        llr_in_tmp[14][39]  = llr_new[14][39];
        llr_in_tmp[14][40]  = llr_new[14][40];
        llr_in_tmp[14][41]  = llr_new[14][41];
    end
 
    2:begin 
        llr_in_tmp[14][0]  = llr_new[14][0];
        llr_in_tmp[14][1]  = llr_new[14][1];
        llr_in_tmp[14][2]  = llr_new[14][2];
        llr_in_tmp[14][3]  = llr_new[14][3];
        llr_in_tmp[14][4]  = llr_new[14][4];
        llr_in_tmp[14][5]  = llr_new[14][5];
        llr_in_tmp[14][6]  = llr_new[14][6];
        llr_in_tmp[14][7]  = llr_new[14][7];
        llr_in_tmp[14][8]  = llr_new[14][8];
        llr_in_tmp[14][9]  = llr_new[14][9];
        llr_in_tmp[14][10]  = llr_new[14][10];
        llr_in_tmp[14][11]  = llr_new[14][11];
        llr_in_tmp[14][12]  = llr_new[14][12];
        llr_in_tmp[14][13]  = llr_new[14][13];
        llr_in_tmp[14][14]  = llr_new[14][14];
        llr_in_tmp[14][15]  = llr_new[14][15];
        llr_in_tmp[14][16]  = llr_new[14][16];
        llr_in_tmp[14][17]  = llr_new[14][17];
        llr_in_tmp[14][18]  = llr_new[14][18];
        llr_in_tmp[14][19]  = llr_new[14][19];
        llr_in_tmp[14][20]  = llr_new[14][20];
        llr_in_tmp[14][21]  = llr_new[14][21];
        llr_in_tmp[14][22]  = llr_new[14][22];
        llr_in_tmp[14][23]  = llr_new[14][23];
        llr_in_tmp[14][24]  = llr_new[14][24];
        llr_in_tmp[14][25]  = llr_new[14][25];
        llr_in_tmp[14][26]  = llr_new[14][26];
        llr_in_tmp[14][27]  = llr_new[14][27];
        llr_in_tmp[14][28]  = llr_new[14][28];
        llr_in_tmp[14][29]  = llr_new[14][29];
        llr_in_tmp[14][30]  = llr_new[14][30];
        llr_in_tmp[14][31]  = llr_new[14][31];
        llr_in_tmp[14][32]  = llr_new[14][32];
        llr_in_tmp[14][33]  = llr_new[14][33];
        llr_in_tmp[14][34]  = llr_new[14][34];
        llr_in_tmp[14][35]  = llr_new[14][35];
        llr_in_tmp[14][36]  = llr_new[14][36];
        llr_in_tmp[14][37]  = llr_new[14][37];
        llr_in_tmp[14][38]  = llr_new[14][38];
        llr_in_tmp[14][39]  = llr_new[14][39];
        llr_in_tmp[14][40]  = llr_new[14][40];
        llr_in_tmp[14][41]  = llr_new[14][41];
    end
 
    3:begin 
        llr_in_tmp[14][0]  = llr_new[14][0];
        llr_in_tmp[14][1]  = llr_new[14][1];
        llr_in_tmp[14][2]  = llr_new[14][2];
        llr_in_tmp[14][3]  = llr_new[14][3];
        llr_in_tmp[14][4]  = llr_new[14][4];
        llr_in_tmp[14][5]  = llr_new[14][5];
        llr_in_tmp[14][6]  = llr_new[14][6];
        llr_in_tmp[14][7]  = llr_new[14][7];
        llr_in_tmp[14][8]  = llr_new[14][8];
        llr_in_tmp[14][9]  = llr_new[14][9];
        llr_in_tmp[14][10]  = llr_new[14][10];
        llr_in_tmp[14][11]  = llr_new[14][11];
        llr_in_tmp[14][12]  = llr_new[14][12];
        llr_in_tmp[14][13]  = llr_new[14][13];
        llr_in_tmp[14][14]  = llr_new[14][14];
        llr_in_tmp[14][15]  = llr_new[14][15];
        llr_in_tmp[14][16]  = llr_new[14][16];
        llr_in_tmp[14][17]  = llr_new[14][17];
        llr_in_tmp[14][18]  = llr_new[14][18];
        llr_in_tmp[14][19]  = llr_new[14][19];
        llr_in_tmp[14][20]  = llr_new[14][20];
        llr_in_tmp[14][21]  = llr_new[14][21];
        llr_in_tmp[14][22]  = llr_new[14][22];
        llr_in_tmp[14][23]  = llr_new[14][23];
        llr_in_tmp[14][24]  = llr_new[14][24];
        llr_in_tmp[14][25]  = llr_new[14][25];
        llr_in_tmp[14][26]  = llr_new[14][26];
        llr_in_tmp[14][27]  = llr_new[14][27];
        llr_in_tmp[14][28]  = llr_new[14][28];
        llr_in_tmp[14][29]  = llr_new[14][29];
        llr_in_tmp[14][30]  = llr_new[14][30];
        llr_in_tmp[14][31]  = llr_new[14][31];
        llr_in_tmp[14][32]  = llr_new[14][32];
        llr_in_tmp[14][33]  = llr_new[14][33];
        llr_in_tmp[14][34]  = llr_new[14][34];
        llr_in_tmp[14][35]  = llr_new[14][35];
        llr_in_tmp[14][36]  = llr_new[14][36];
        llr_in_tmp[14][37]  = llr_new[14][37];
        llr_in_tmp[14][38]  = llr_new[14][38];
        llr_in_tmp[14][39]  = llr_new[14][39];
        llr_in_tmp[14][40]  = llr_new[14][40];
        llr_in_tmp[14][41]  = llr_new[14][41];
    end
 
    4:begin 
        llr_in_tmp[14][0]  = llr_new[14][0];
        llr_in_tmp[14][1]  = llr_new[14][1];
        llr_in_tmp[14][2]  = llr_new[14][2];
        llr_in_tmp[14][3]  = llr_new[14][3];
        llr_in_tmp[14][4]  = llr_new[14][4];
        llr_in_tmp[14][5]  = llr_new[14][5];
        llr_in_tmp[14][6]  = llr_new[14][6];
        llr_in_tmp[14][7]  = llr_new[14][7];
        llr_in_tmp[14][8]  = llr_new[14][8];
        llr_in_tmp[14][9]  = llr_new[14][9];
        llr_in_tmp[14][10]  = llr_new[14][10];
        llr_in_tmp[14][11]  = llr_new[14][11];
        llr_in_tmp[14][12]  = llr_new[14][12];
        llr_in_tmp[14][13]  = llr_new[14][13];
        llr_in_tmp[14][14]  = llr_new[14][14];
        llr_in_tmp[14][15]  = llr_new[14][15];
        llr_in_tmp[14][16]  = llr_new[14][16];
        llr_in_tmp[14][17]  = llr_new[14][17];
        llr_in_tmp[14][18]  = llr_new[14][18];
        llr_in_tmp[14][19]  = llr_new[14][19];
        llr_in_tmp[14][20]  = llr_new[14][20];
        llr_in_tmp[14][21]  = llr_new[14][21];
        llr_in_tmp[14][22]  = llr_new[14][22];
        llr_in_tmp[14][23]  = llr_new[14][23];
        llr_in_tmp[14][24]  = llr_new[14][24];
        llr_in_tmp[14][25]  = llr_new[14][25];
        llr_in_tmp[14][26]  = llr_new[14][26];
        llr_in_tmp[14][27]  = llr_new[14][27];
        llr_in_tmp[14][28]  = llr_new[14][28];
        llr_in_tmp[14][29]  = llr_new[14][29];
        llr_in_tmp[14][30]  = llr_new[14][30];
        llr_in_tmp[14][31]  = llr_new[14][31];
        llr_in_tmp[14][32]  = llr_new[14][32];
        llr_in_tmp[14][33]  = llr_new[14][33];
        llr_in_tmp[14][34]  = llr_new[14][34];
        llr_in_tmp[14][35]  = llr_new[14][35];
        llr_in_tmp[14][36]  = llr_new[14][36];
        llr_in_tmp[14][37]  = llr_new[14][37];
        llr_in_tmp[14][38]  = llr_new[14][38];
        llr_in_tmp[14][39]  = llr_new[14][39];
        llr_in_tmp[14][40]  = llr_new[14][40];
        llr_in_tmp[14][41]  = llr_new[14][41];
    end
 
    5:begin 
        llr_in_tmp[14][0]  = llr_new[14][0];
        llr_in_tmp[14][1]  = llr_new[14][1];
        llr_in_tmp[14][2]  = llr_new[14][2];
        llr_in_tmp[14][3]  = llr_new[14][3];
        llr_in_tmp[14][4]  = llr_new[14][4];
        llr_in_tmp[14][5]  = llr_new[14][5];
        llr_in_tmp[14][6]  = llr_new[14][6];
        llr_in_tmp[14][7]  = llr_new[14][7];
        llr_in_tmp[14][8]  = llr_new[14][8];
        llr_in_tmp[14][9]  = llr_new[14][9];
        llr_in_tmp[14][10]  = llr_new[14][10];
        llr_in_tmp[14][11]  = llr_new[14][11];
        llr_in_tmp[14][12]  = llr_new[14][12];
        llr_in_tmp[14][13]  = llr_new[14][13];
        llr_in_tmp[14][14]  = llr_new[14][14];
        llr_in_tmp[14][15]  = llr_new[14][15];
        llr_in_tmp[14][16]  = llr_new[14][16];
        llr_in_tmp[14][17]  = llr_new[14][17];
        llr_in_tmp[14][18]  = llr_new[14][18];
        llr_in_tmp[14][19]  = llr_new[14][19];
        llr_in_tmp[14][20]  = llr_new[14][20];
        llr_in_tmp[14][21]  = llr_new[14][21];
        llr_in_tmp[14][22]  = llr_new[14][22];
        llr_in_tmp[14][23]  = llr_new[14][23];
        llr_in_tmp[14][24]  = llr_new[14][24];
        llr_in_tmp[14][25]  = llr_new[14][25];
        llr_in_tmp[14][26]  = llr_new[14][26];
        llr_in_tmp[14][27]  = llr_new[14][27];
        llr_in_tmp[14][28]  = llr_new[14][28];
        llr_in_tmp[14][29]  = llr_new[14][29];
        llr_in_tmp[14][30]  = llr_new[14][30];
        llr_in_tmp[14][31]  = llr_new[14][31];
        llr_in_tmp[14][32]  = llr_new[14][32];
        llr_in_tmp[14][33]  = llr_new[14][33];
        llr_in_tmp[14][34]  = llr_new[14][34];
        llr_in_tmp[14][35]  = llr_new[14][35];
        llr_in_tmp[14][36]  = llr_new[14][36];
        llr_in_tmp[14][37]  = llr_new[14][37];
        llr_in_tmp[14][38]  = llr_new[14][38];
        llr_in_tmp[14][39]  = llr_new[14][39];
        llr_in_tmp[14][40]  = llr_new[14][40];
        llr_in_tmp[14][41]  = llr_new[14][41];
    end
 
    6:begin 
        llr_in_tmp[14][0]  = llr_new[14][13];
        llr_in_tmp[14][1]  = llr_new[14][14];
        llr_in_tmp[14][2]  = llr_new[14][15];
        llr_in_tmp[14][3]  = llr_new[14][16];
        llr_in_tmp[14][4]  = llr_new[14][17];
        llr_in_tmp[14][5]  = llr_new[14][18];
        llr_in_tmp[14][6]  = llr_new[14][19];
        llr_in_tmp[14][7]  = llr_new[14][20];
        llr_in_tmp[14][8]  = llr_new[14][21];
        llr_in_tmp[14][9]  = llr_new[14][22];
        llr_in_tmp[14][10]  = llr_new[14][23];
        llr_in_tmp[14][11]  = llr_new[14][24];
        llr_in_tmp[14][12]  = llr_new[14][25];
        llr_in_tmp[14][13]  = llr_new[14][26];
        llr_in_tmp[14][14]  = llr_new[14][27];
        llr_in_tmp[14][15]  = llr_new[14][28];
        llr_in_tmp[14][16]  = llr_new[14][29];
        llr_in_tmp[14][17]  = llr_new[14][30];
        llr_in_tmp[14][18]  = llr_new[14][31];
        llr_in_tmp[14][19]  = llr_new[14][32];
        llr_in_tmp[14][20]  = llr_new[14][33];
        llr_in_tmp[14][21]  = llr_new[14][34];
        llr_in_tmp[14][22]  = llr_new[14][35];
        llr_in_tmp[14][23]  = llr_new[14][36];
        llr_in_tmp[14][24]  = llr_new[14][37];
        llr_in_tmp[14][25]  = llr_new[14][38];
        llr_in_tmp[14][26]  = llr_new[14][39];
        llr_in_tmp[14][27]  = llr_new[14][40];
        llr_in_tmp[14][28]  = llr_new[14][41];
        llr_in_tmp[14][29]  = llr_new[14][0];
        llr_in_tmp[14][30]  = llr_new[14][1];
        llr_in_tmp[14][31]  = llr_new[14][2];
        llr_in_tmp[14][32]  = llr_new[14][3];
        llr_in_tmp[14][33]  = llr_new[14][4];
        llr_in_tmp[14][34]  = llr_new[14][5];
        llr_in_tmp[14][35]  = llr_new[14][6];
        llr_in_tmp[14][36]  = llr_new[14][7];
        llr_in_tmp[14][37]  = llr_new[14][8];
        llr_in_tmp[14][38]  = llr_new[14][9];
        llr_in_tmp[14][39]  = llr_new[14][10];
        llr_in_tmp[14][40]  = llr_new[14][11];
        llr_in_tmp[14][41]  = llr_new[14][12];
    end
 
    7:begin 
        llr_in_tmp[14][0]  = llr_new[14][22];
        llr_in_tmp[14][1]  = llr_new[14][23];
        llr_in_tmp[14][2]  = llr_new[14][24];
        llr_in_tmp[14][3]  = llr_new[14][25];
        llr_in_tmp[14][4]  = llr_new[14][26];
        llr_in_tmp[14][5]  = llr_new[14][27];
        llr_in_tmp[14][6]  = llr_new[14][28];
        llr_in_tmp[14][7]  = llr_new[14][29];
        llr_in_tmp[14][8]  = llr_new[14][30];
        llr_in_tmp[14][9]  = llr_new[14][31];
        llr_in_tmp[14][10]  = llr_new[14][32];
        llr_in_tmp[14][11]  = llr_new[14][33];
        llr_in_tmp[14][12]  = llr_new[14][34];
        llr_in_tmp[14][13]  = llr_new[14][35];
        llr_in_tmp[14][14]  = llr_new[14][36];
        llr_in_tmp[14][15]  = llr_new[14][37];
        llr_in_tmp[14][16]  = llr_new[14][38];
        llr_in_tmp[14][17]  = llr_new[14][39];
        llr_in_tmp[14][18]  = llr_new[14][40];
        llr_in_tmp[14][19]  = llr_new[14][41];
        llr_in_tmp[14][20]  = llr_new[14][0];
        llr_in_tmp[14][21]  = llr_new[14][1];
        llr_in_tmp[14][22]  = llr_new[14][2];
        llr_in_tmp[14][23]  = llr_new[14][3];
        llr_in_tmp[14][24]  = llr_new[14][4];
        llr_in_tmp[14][25]  = llr_new[14][5];
        llr_in_tmp[14][26]  = llr_new[14][6];
        llr_in_tmp[14][27]  = llr_new[14][7];
        llr_in_tmp[14][28]  = llr_new[14][8];
        llr_in_tmp[14][29]  = llr_new[14][9];
        llr_in_tmp[14][30]  = llr_new[14][10];
        llr_in_tmp[14][31]  = llr_new[14][11];
        llr_in_tmp[14][32]  = llr_new[14][12];
        llr_in_tmp[14][33]  = llr_new[14][13];
        llr_in_tmp[14][34]  = llr_new[14][14];
        llr_in_tmp[14][35]  = llr_new[14][15];
        llr_in_tmp[14][36]  = llr_new[14][16];
        llr_in_tmp[14][37]  = llr_new[14][17];
        llr_in_tmp[14][38]  = llr_new[14][18];
        llr_in_tmp[14][39]  = llr_new[14][19];
        llr_in_tmp[14][40]  = llr_new[14][20];
        llr_in_tmp[14][41]  = llr_new[14][21];
    end
 
endcase
end

if (chk_n_input_valid) begin
case (curr_layer)
    0:begin 
        llr_in_tmp[15][0]  = llr_new[15][0];
        llr_in_tmp[15][1]  = llr_new[15][1];
        llr_in_tmp[15][2]  = llr_new[15][2];
        llr_in_tmp[15][3]  = llr_new[15][3];
        llr_in_tmp[15][4]  = llr_new[15][4];
        llr_in_tmp[15][5]  = llr_new[15][5];
        llr_in_tmp[15][6]  = llr_new[15][6];
        llr_in_tmp[15][7]  = llr_new[15][7];
        llr_in_tmp[15][8]  = llr_new[15][8];
        llr_in_tmp[15][9]  = llr_new[15][9];
        llr_in_tmp[15][10]  = llr_new[15][10];
        llr_in_tmp[15][11]  = llr_new[15][11];
        llr_in_tmp[15][12]  = llr_new[15][12];
        llr_in_tmp[15][13]  = llr_new[15][13];
        llr_in_tmp[15][14]  = llr_new[15][14];
        llr_in_tmp[15][15]  = llr_new[15][15];
        llr_in_tmp[15][16]  = llr_new[15][16];
        llr_in_tmp[15][17]  = llr_new[15][17];
        llr_in_tmp[15][18]  = llr_new[15][18];
        llr_in_tmp[15][19]  = llr_new[15][19];
        llr_in_tmp[15][20]  = llr_new[15][20];
        llr_in_tmp[15][21]  = llr_new[15][21];
        llr_in_tmp[15][22]  = llr_new[15][22];
        llr_in_tmp[15][23]  = llr_new[15][23];
        llr_in_tmp[15][24]  = llr_new[15][24];
        llr_in_tmp[15][25]  = llr_new[15][25];
        llr_in_tmp[15][26]  = llr_new[15][26];
        llr_in_tmp[15][27]  = llr_new[15][27];
        llr_in_tmp[15][28]  = llr_new[15][28];
        llr_in_tmp[15][29]  = llr_new[15][29];
        llr_in_tmp[15][30]  = llr_new[15][30];
        llr_in_tmp[15][31]  = llr_new[15][31];
        llr_in_tmp[15][32]  = llr_new[15][32];
        llr_in_tmp[15][33]  = llr_new[15][33];
        llr_in_tmp[15][34]  = llr_new[15][34];
        llr_in_tmp[15][35]  = llr_new[15][35];
        llr_in_tmp[15][36]  = llr_new[15][36];
        llr_in_tmp[15][37]  = llr_new[15][37];
        llr_in_tmp[15][38]  = llr_new[15][38];
        llr_in_tmp[15][39]  = llr_new[15][39];
        llr_in_tmp[15][40]  = llr_new[15][40];
        llr_in_tmp[15][41]  = llr_new[15][41];
    end
 
    1:begin 
        llr_in_tmp[15][0]  = llr_new[15][0];
        llr_in_tmp[15][1]  = llr_new[15][1];
        llr_in_tmp[15][2]  = llr_new[15][2];
        llr_in_tmp[15][3]  = llr_new[15][3];
        llr_in_tmp[15][4]  = llr_new[15][4];
        llr_in_tmp[15][5]  = llr_new[15][5];
        llr_in_tmp[15][6]  = llr_new[15][6];
        llr_in_tmp[15][7]  = llr_new[15][7];
        llr_in_tmp[15][8]  = llr_new[15][8];
        llr_in_tmp[15][9]  = llr_new[15][9];
        llr_in_tmp[15][10]  = llr_new[15][10];
        llr_in_tmp[15][11]  = llr_new[15][11];
        llr_in_tmp[15][12]  = llr_new[15][12];
        llr_in_tmp[15][13]  = llr_new[15][13];
        llr_in_tmp[15][14]  = llr_new[15][14];
        llr_in_tmp[15][15]  = llr_new[15][15];
        llr_in_tmp[15][16]  = llr_new[15][16];
        llr_in_tmp[15][17]  = llr_new[15][17];
        llr_in_tmp[15][18]  = llr_new[15][18];
        llr_in_tmp[15][19]  = llr_new[15][19];
        llr_in_tmp[15][20]  = llr_new[15][20];
        llr_in_tmp[15][21]  = llr_new[15][21];
        llr_in_tmp[15][22]  = llr_new[15][22];
        llr_in_tmp[15][23]  = llr_new[15][23];
        llr_in_tmp[15][24]  = llr_new[15][24];
        llr_in_tmp[15][25]  = llr_new[15][25];
        llr_in_tmp[15][26]  = llr_new[15][26];
        llr_in_tmp[15][27]  = llr_new[15][27];
        llr_in_tmp[15][28]  = llr_new[15][28];
        llr_in_tmp[15][29]  = llr_new[15][29];
        llr_in_tmp[15][30]  = llr_new[15][30];
        llr_in_tmp[15][31]  = llr_new[15][31];
        llr_in_tmp[15][32]  = llr_new[15][32];
        llr_in_tmp[15][33]  = llr_new[15][33];
        llr_in_tmp[15][34]  = llr_new[15][34];
        llr_in_tmp[15][35]  = llr_new[15][35];
        llr_in_tmp[15][36]  = llr_new[15][36];
        llr_in_tmp[15][37]  = llr_new[15][37];
        llr_in_tmp[15][38]  = llr_new[15][38];
        llr_in_tmp[15][39]  = llr_new[15][39];
        llr_in_tmp[15][40]  = llr_new[15][40];
        llr_in_tmp[15][41]  = llr_new[15][41];
    end
 
    2:begin 
        llr_in_tmp[15][0]  = llr_new[15][0];
        llr_in_tmp[15][1]  = llr_new[15][1];
        llr_in_tmp[15][2]  = llr_new[15][2];
        llr_in_tmp[15][3]  = llr_new[15][3];
        llr_in_tmp[15][4]  = llr_new[15][4];
        llr_in_tmp[15][5]  = llr_new[15][5];
        llr_in_tmp[15][6]  = llr_new[15][6];
        llr_in_tmp[15][7]  = llr_new[15][7];
        llr_in_tmp[15][8]  = llr_new[15][8];
        llr_in_tmp[15][9]  = llr_new[15][9];
        llr_in_tmp[15][10]  = llr_new[15][10];
        llr_in_tmp[15][11]  = llr_new[15][11];
        llr_in_tmp[15][12]  = llr_new[15][12];
        llr_in_tmp[15][13]  = llr_new[15][13];
        llr_in_tmp[15][14]  = llr_new[15][14];
        llr_in_tmp[15][15]  = llr_new[15][15];
        llr_in_tmp[15][16]  = llr_new[15][16];
        llr_in_tmp[15][17]  = llr_new[15][17];
        llr_in_tmp[15][18]  = llr_new[15][18];
        llr_in_tmp[15][19]  = llr_new[15][19];
        llr_in_tmp[15][20]  = llr_new[15][20];
        llr_in_tmp[15][21]  = llr_new[15][21];
        llr_in_tmp[15][22]  = llr_new[15][22];
        llr_in_tmp[15][23]  = llr_new[15][23];
        llr_in_tmp[15][24]  = llr_new[15][24];
        llr_in_tmp[15][25]  = llr_new[15][25];
        llr_in_tmp[15][26]  = llr_new[15][26];
        llr_in_tmp[15][27]  = llr_new[15][27];
        llr_in_tmp[15][28]  = llr_new[15][28];
        llr_in_tmp[15][29]  = llr_new[15][29];
        llr_in_tmp[15][30]  = llr_new[15][30];
        llr_in_tmp[15][31]  = llr_new[15][31];
        llr_in_tmp[15][32]  = llr_new[15][32];
        llr_in_tmp[15][33]  = llr_new[15][33];
        llr_in_tmp[15][34]  = llr_new[15][34];
        llr_in_tmp[15][35]  = llr_new[15][35];
        llr_in_tmp[15][36]  = llr_new[15][36];
        llr_in_tmp[15][37]  = llr_new[15][37];
        llr_in_tmp[15][38]  = llr_new[15][38];
        llr_in_tmp[15][39]  = llr_new[15][39];
        llr_in_tmp[15][40]  = llr_new[15][40];
        llr_in_tmp[15][41]  = llr_new[15][41];
    end
 
    3:begin 
        llr_in_tmp[15][0]  = llr_new[15][0];
        llr_in_tmp[15][1]  = llr_new[15][1];
        llr_in_tmp[15][2]  = llr_new[15][2];
        llr_in_tmp[15][3]  = llr_new[15][3];
        llr_in_tmp[15][4]  = llr_new[15][4];
        llr_in_tmp[15][5]  = llr_new[15][5];
        llr_in_tmp[15][6]  = llr_new[15][6];
        llr_in_tmp[15][7]  = llr_new[15][7];
        llr_in_tmp[15][8]  = llr_new[15][8];
        llr_in_tmp[15][9]  = llr_new[15][9];
        llr_in_tmp[15][10]  = llr_new[15][10];
        llr_in_tmp[15][11]  = llr_new[15][11];
        llr_in_tmp[15][12]  = llr_new[15][12];
        llr_in_tmp[15][13]  = llr_new[15][13];
        llr_in_tmp[15][14]  = llr_new[15][14];
        llr_in_tmp[15][15]  = llr_new[15][15];
        llr_in_tmp[15][16]  = llr_new[15][16];
        llr_in_tmp[15][17]  = llr_new[15][17];
        llr_in_tmp[15][18]  = llr_new[15][18];
        llr_in_tmp[15][19]  = llr_new[15][19];
        llr_in_tmp[15][20]  = llr_new[15][20];
        llr_in_tmp[15][21]  = llr_new[15][21];
        llr_in_tmp[15][22]  = llr_new[15][22];
        llr_in_tmp[15][23]  = llr_new[15][23];
        llr_in_tmp[15][24]  = llr_new[15][24];
        llr_in_tmp[15][25]  = llr_new[15][25];
        llr_in_tmp[15][26]  = llr_new[15][26];
        llr_in_tmp[15][27]  = llr_new[15][27];
        llr_in_tmp[15][28]  = llr_new[15][28];
        llr_in_tmp[15][29]  = llr_new[15][29];
        llr_in_tmp[15][30]  = llr_new[15][30];
        llr_in_tmp[15][31]  = llr_new[15][31];
        llr_in_tmp[15][32]  = llr_new[15][32];
        llr_in_tmp[15][33]  = llr_new[15][33];
        llr_in_tmp[15][34]  = llr_new[15][34];
        llr_in_tmp[15][35]  = llr_new[15][35];
        llr_in_tmp[15][36]  = llr_new[15][36];
        llr_in_tmp[15][37]  = llr_new[15][37];
        llr_in_tmp[15][38]  = llr_new[15][38];
        llr_in_tmp[15][39]  = llr_new[15][39];
        llr_in_tmp[15][40]  = llr_new[15][40];
        llr_in_tmp[15][41]  = llr_new[15][41];
    end
 
    4:begin 
        llr_in_tmp[15][0]  = llr_new[15][0];
        llr_in_tmp[15][1]  = llr_new[15][1];
        llr_in_tmp[15][2]  = llr_new[15][2];
        llr_in_tmp[15][3]  = llr_new[15][3];
        llr_in_tmp[15][4]  = llr_new[15][4];
        llr_in_tmp[15][5]  = llr_new[15][5];
        llr_in_tmp[15][6]  = llr_new[15][6];
        llr_in_tmp[15][7]  = llr_new[15][7];
        llr_in_tmp[15][8]  = llr_new[15][8];
        llr_in_tmp[15][9]  = llr_new[15][9];
        llr_in_tmp[15][10]  = llr_new[15][10];
        llr_in_tmp[15][11]  = llr_new[15][11];
        llr_in_tmp[15][12]  = llr_new[15][12];
        llr_in_tmp[15][13]  = llr_new[15][13];
        llr_in_tmp[15][14]  = llr_new[15][14];
        llr_in_tmp[15][15]  = llr_new[15][15];
        llr_in_tmp[15][16]  = llr_new[15][16];
        llr_in_tmp[15][17]  = llr_new[15][17];
        llr_in_tmp[15][18]  = llr_new[15][18];
        llr_in_tmp[15][19]  = llr_new[15][19];
        llr_in_tmp[15][20]  = llr_new[15][20];
        llr_in_tmp[15][21]  = llr_new[15][21];
        llr_in_tmp[15][22]  = llr_new[15][22];
        llr_in_tmp[15][23]  = llr_new[15][23];
        llr_in_tmp[15][24]  = llr_new[15][24];
        llr_in_tmp[15][25]  = llr_new[15][25];
        llr_in_tmp[15][26]  = llr_new[15][26];
        llr_in_tmp[15][27]  = llr_new[15][27];
        llr_in_tmp[15][28]  = llr_new[15][28];
        llr_in_tmp[15][29]  = llr_new[15][29];
        llr_in_tmp[15][30]  = llr_new[15][30];
        llr_in_tmp[15][31]  = llr_new[15][31];
        llr_in_tmp[15][32]  = llr_new[15][32];
        llr_in_tmp[15][33]  = llr_new[15][33];
        llr_in_tmp[15][34]  = llr_new[15][34];
        llr_in_tmp[15][35]  = llr_new[15][35];
        llr_in_tmp[15][36]  = llr_new[15][36];
        llr_in_tmp[15][37]  = llr_new[15][37];
        llr_in_tmp[15][38]  = llr_new[15][38];
        llr_in_tmp[15][39]  = llr_new[15][39];
        llr_in_tmp[15][40]  = llr_new[15][40];
        llr_in_tmp[15][41]  = llr_new[15][41];
    end
 
    5:begin 
        llr_in_tmp[15][0]  = llr_new[15][0];
        llr_in_tmp[15][1]  = llr_new[15][1];
        llr_in_tmp[15][2]  = llr_new[15][2];
        llr_in_tmp[15][3]  = llr_new[15][3];
        llr_in_tmp[15][4]  = llr_new[15][4];
        llr_in_tmp[15][5]  = llr_new[15][5];
        llr_in_tmp[15][6]  = llr_new[15][6];
        llr_in_tmp[15][7]  = llr_new[15][7];
        llr_in_tmp[15][8]  = llr_new[15][8];
        llr_in_tmp[15][9]  = llr_new[15][9];
        llr_in_tmp[15][10]  = llr_new[15][10];
        llr_in_tmp[15][11]  = llr_new[15][11];
        llr_in_tmp[15][12]  = llr_new[15][12];
        llr_in_tmp[15][13]  = llr_new[15][13];
        llr_in_tmp[15][14]  = llr_new[15][14];
        llr_in_tmp[15][15]  = llr_new[15][15];
        llr_in_tmp[15][16]  = llr_new[15][16];
        llr_in_tmp[15][17]  = llr_new[15][17];
        llr_in_tmp[15][18]  = llr_new[15][18];
        llr_in_tmp[15][19]  = llr_new[15][19];
        llr_in_tmp[15][20]  = llr_new[15][20];
        llr_in_tmp[15][21]  = llr_new[15][21];
        llr_in_tmp[15][22]  = llr_new[15][22];
        llr_in_tmp[15][23]  = llr_new[15][23];
        llr_in_tmp[15][24]  = llr_new[15][24];
        llr_in_tmp[15][25]  = llr_new[15][25];
        llr_in_tmp[15][26]  = llr_new[15][26];
        llr_in_tmp[15][27]  = llr_new[15][27];
        llr_in_tmp[15][28]  = llr_new[15][28];
        llr_in_tmp[15][29]  = llr_new[15][29];
        llr_in_tmp[15][30]  = llr_new[15][30];
        llr_in_tmp[15][31]  = llr_new[15][31];
        llr_in_tmp[15][32]  = llr_new[15][32];
        llr_in_tmp[15][33]  = llr_new[15][33];
        llr_in_tmp[15][34]  = llr_new[15][34];
        llr_in_tmp[15][35]  = llr_new[15][35];
        llr_in_tmp[15][36]  = llr_new[15][36];
        llr_in_tmp[15][37]  = llr_new[15][37];
        llr_in_tmp[15][38]  = llr_new[15][38];
        llr_in_tmp[15][39]  = llr_new[15][39];
        llr_in_tmp[15][40]  = llr_new[15][40];
        llr_in_tmp[15][41]  = llr_new[15][41];
    end
 
    6:begin 
        llr_in_tmp[15][0]  = llr_new[15][0];
        llr_in_tmp[15][1]  = llr_new[15][1];
        llr_in_tmp[15][2]  = llr_new[15][2];
        llr_in_tmp[15][3]  = llr_new[15][3];
        llr_in_tmp[15][4]  = llr_new[15][4];
        llr_in_tmp[15][5]  = llr_new[15][5];
        llr_in_tmp[15][6]  = llr_new[15][6];
        llr_in_tmp[15][7]  = llr_new[15][7];
        llr_in_tmp[15][8]  = llr_new[15][8];
        llr_in_tmp[15][9]  = llr_new[15][9];
        llr_in_tmp[15][10]  = llr_new[15][10];
        llr_in_tmp[15][11]  = llr_new[15][11];
        llr_in_tmp[15][12]  = llr_new[15][12];
        llr_in_tmp[15][13]  = llr_new[15][13];
        llr_in_tmp[15][14]  = llr_new[15][14];
        llr_in_tmp[15][15]  = llr_new[15][15];
        llr_in_tmp[15][16]  = llr_new[15][16];
        llr_in_tmp[15][17]  = llr_new[15][17];
        llr_in_tmp[15][18]  = llr_new[15][18];
        llr_in_tmp[15][19]  = llr_new[15][19];
        llr_in_tmp[15][20]  = llr_new[15][20];
        llr_in_tmp[15][21]  = llr_new[15][21];
        llr_in_tmp[15][22]  = llr_new[15][22];
        llr_in_tmp[15][23]  = llr_new[15][23];
        llr_in_tmp[15][24]  = llr_new[15][24];
        llr_in_tmp[15][25]  = llr_new[15][25];
        llr_in_tmp[15][26]  = llr_new[15][26];
        llr_in_tmp[15][27]  = llr_new[15][27];
        llr_in_tmp[15][28]  = llr_new[15][28];
        llr_in_tmp[15][29]  = llr_new[15][29];
        llr_in_tmp[15][30]  = llr_new[15][30];
        llr_in_tmp[15][31]  = llr_new[15][31];
        llr_in_tmp[15][32]  = llr_new[15][32];
        llr_in_tmp[15][33]  = llr_new[15][33];
        llr_in_tmp[15][34]  = llr_new[15][34];
        llr_in_tmp[15][35]  = llr_new[15][35];
        llr_in_tmp[15][36]  = llr_new[15][36];
        llr_in_tmp[15][37]  = llr_new[15][37];
        llr_in_tmp[15][38]  = llr_new[15][38];
        llr_in_tmp[15][39]  = llr_new[15][39];
        llr_in_tmp[15][40]  = llr_new[15][40];
        llr_in_tmp[15][41]  = llr_new[15][41];
    end
 
    7:begin 
        llr_in_tmp[15][0]  = llr_new[15][24];
        llr_in_tmp[15][1]  = llr_new[15][25];
        llr_in_tmp[15][2]  = llr_new[15][26];
        llr_in_tmp[15][3]  = llr_new[15][27];
        llr_in_tmp[15][4]  = llr_new[15][28];
        llr_in_tmp[15][5]  = llr_new[15][29];
        llr_in_tmp[15][6]  = llr_new[15][30];
        llr_in_tmp[15][7]  = llr_new[15][31];
        llr_in_tmp[15][8]  = llr_new[15][32];
        llr_in_tmp[15][9]  = llr_new[15][33];
        llr_in_tmp[15][10]  = llr_new[15][34];
        llr_in_tmp[15][11]  = llr_new[15][35];
        llr_in_tmp[15][12]  = llr_new[15][36];
        llr_in_tmp[15][13]  = llr_new[15][37];
        llr_in_tmp[15][14]  = llr_new[15][38];
        llr_in_tmp[15][15]  = llr_new[15][39];
        llr_in_tmp[15][16]  = llr_new[15][40];
        llr_in_tmp[15][17]  = llr_new[15][41];
        llr_in_tmp[15][18]  = llr_new[15][0];
        llr_in_tmp[15][19]  = llr_new[15][1];
        llr_in_tmp[15][20]  = llr_new[15][2];
        llr_in_tmp[15][21]  = llr_new[15][3];
        llr_in_tmp[15][22]  = llr_new[15][4];
        llr_in_tmp[15][23]  = llr_new[15][5];
        llr_in_tmp[15][24]  = llr_new[15][6];
        llr_in_tmp[15][25]  = llr_new[15][7];
        llr_in_tmp[15][26]  = llr_new[15][8];
        llr_in_tmp[15][27]  = llr_new[15][9];
        llr_in_tmp[15][28]  = llr_new[15][10];
        llr_in_tmp[15][29]  = llr_new[15][11];
        llr_in_tmp[15][30]  = llr_new[15][12];
        llr_in_tmp[15][31]  = llr_new[15][13];
        llr_in_tmp[15][32]  = llr_new[15][14];
        llr_in_tmp[15][33]  = llr_new[15][15];
        llr_in_tmp[15][34]  = llr_new[15][16];
        llr_in_tmp[15][35]  = llr_new[15][17];
        llr_in_tmp[15][36]  = llr_new[15][18];
        llr_in_tmp[15][37]  = llr_new[15][19];
        llr_in_tmp[15][38]  = llr_new[15][20];
        llr_in_tmp[15][39]  = llr_new[15][21];
        llr_in_tmp[15][40]  = llr_new[15][22];
        llr_in_tmp[15][41]  = llr_new[15][23];
    end
 
endcase
end

end
